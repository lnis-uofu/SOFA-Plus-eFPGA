//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Formal Top-level netlist of Design: counter
//	 removed 
//	Organization: University of Utah
//	 removed 
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
// `default_nettype wire

module counter_top_formal_verification_random_tb;
// ----- Default clock port is added here since benchmark does not contain one -------
	reg [0:0] clk;

// ----- Shared inputs -------
	reg [0:0] resetb;

// ----- FPGA fabric outputs -------
	wire [0:0] out_result_0__gfpga;
	wire [0:0] out_result_1__gfpga;
	wire [0:0] out_result_2__gfpga;
	wire [0:0] out_result_3__gfpga;
	wire [0:0] out_result_4__gfpga;
	wire [0:0] out_result_5__gfpga;
	wire [0:0] out_result_6__gfpga;
	wire [0:0] out_result_7__gfpga;
	wire [0:0] out_result_8__gfpga;
	wire [0:0] out_result_9__gfpga;
	wire [0:0] out_result_10__gfpga;
	wire [0:0] out_result_11__gfpga;
	wire [0:0] out_result_12__gfpga;
	wire [0:0] out_result_13__gfpga;
	wire [0:0] out_result_14__gfpga;
	wire [0:0] out_result_15__gfpga;
	wire [0:0] out_result_16__gfpga;
	wire [0:0] out_result_17__gfpga;
	wire [0:0] out_result_18__gfpga;
	wire [0:0] out_result_19__gfpga;
	wire [0:0] out_result_20__gfpga;
	wire [0:0] out_result_21__gfpga;
	wire [0:0] out_result_22__gfpga;
	wire [0:0] out_result_23__gfpga;
	wire [0:0] out_result_24__gfpga;
	wire [0:0] out_result_25__gfpga;
	wire [0:0] out_result_26__gfpga;
	wire [0:0] out_result_27__gfpga;
	wire [0:0] out_result_28__gfpga;
	wire [0:0] out_result_29__gfpga;
	wire [0:0] out_result_30__gfpga;
	wire [0:0] out_result_31__gfpga;
	wire [0:0] out_result_32__gfpga;
	wire [0:0] out_result_33__gfpga;
	wire [0:0] out_result_34__gfpga;
	wire [0:0] out_result_35__gfpga;
	wire [0:0] out_result_36__gfpga;
	wire [0:0] out_result_37__gfpga;
	wire [0:0] out_result_38__gfpga;
	wire [0:0] out_result_39__gfpga;
	wire [0:0] out_result_40__gfpga;
	wire [0:0] out_result_41__gfpga;
	wire [0:0] out_result_42__gfpga;
	wire [0:0] out_result_43__gfpga;
	wire [0:0] out_result_44__gfpga;
	wire [0:0] out_result_45__gfpga;
	wire [0:0] out_result_46__gfpga;
	wire [0:0] out_result_47__gfpga;
	wire [0:0] out_result_48__gfpga;
	wire [0:0] out_result_49__gfpga;
	wire [0:0] out_result_50__gfpga;
	wire [0:0] out_result_51__gfpga;
	wire [0:0] out_result_52__gfpga;
	wire [0:0] out_result_53__gfpga;
	wire [0:0] out_result_54__gfpga;
	wire [0:0] out_result_55__gfpga;
	wire [0:0] out_result_56__gfpga;
	wire [0:0] out_result_57__gfpga;
	wire [0:0] out_result_58__gfpga;
	wire [0:0] out_result_59__gfpga;
	wire [0:0] out_result_60__gfpga;
	wire [0:0] out_result_61__gfpga;
	wire [0:0] out_result_62__gfpga;
	wire [0:0] out_result_63__gfpga;
	wire [0:0] out_result_64__gfpga;
	wire [0:0] out_result_65__gfpga;
	wire [0:0] out_result_66__gfpga;
	wire [0:0] out_result_67__gfpga;
	wire [0:0] out_result_68__gfpga;
	wire [0:0] out_result_69__gfpga;
	wire [0:0] out_result_70__gfpga;
	wire [0:0] out_result_71__gfpga;
	wire [0:0] out_result_72__gfpga;
	wire [0:0] out_result_73__gfpga;
	wire [0:0] out_result_74__gfpga;
	wire [0:0] out_result_75__gfpga;
	wire [0:0] out_result_76__gfpga;
	wire [0:0] out_result_77__gfpga;
	wire [0:0] out_result_78__gfpga;
	wire [0:0] out_result_79__gfpga;
	wire [0:0] out_result_80__gfpga;
	wire [0:0] out_result_81__gfpga;
	wire [0:0] out_result_82__gfpga;
	wire [0:0] out_result_83__gfpga;
	wire [0:0] out_result_84__gfpga;
	wire [0:0] out_result_85__gfpga;
	wire [0:0] out_result_86__gfpga;
	wire [0:0] out_result_87__gfpga;
	wire [0:0] out_result_88__gfpga;
	wire [0:0] out_result_89__gfpga;
	wire [0:0] out_result_90__gfpga;
	wire [0:0] out_result_91__gfpga;
	wire [0:0] out_result_92__gfpga;
	wire [0:0] out_result_93__gfpga;
	wire [0:0] out_result_94__gfpga;
	wire [0:0] out_result_95__gfpga;
	wire [0:0] out_result_96__gfpga;
	wire [0:0] out_result_97__gfpga;
	wire [0:0] out_result_98__gfpga;
	wire [0:0] out_result_99__gfpga;
	wire [0:0] out_result_100__gfpga;
	wire [0:0] out_result_101__gfpga;
	wire [0:0] out_result_102__gfpga;
	wire [0:0] out_result_103__gfpga;
	wire [0:0] out_result_104__gfpga;
	wire [0:0] out_result_105__gfpga;
	wire [0:0] out_result_106__gfpga;
	wire [0:0] out_result_107__gfpga;
	wire [0:0] out_result_108__gfpga;
	wire [0:0] out_result_109__gfpga;
	wire [0:0] out_result_110__gfpga;
	wire [0:0] out_result_111__gfpga;
	wire [0:0] out_result_112__gfpga;
	wire [0:0] out_result_113__gfpga;
	wire [0:0] out_result_114__gfpga;
	wire [0:0] out_result_115__gfpga;
	wire [0:0] out_result_116__gfpga;
	wire [0:0] out_result_117__gfpga;
	wire [0:0] out_result_118__gfpga;
	wire [0:0] out_result_119__gfpga;
	wire [0:0] out_result_120__gfpga;
	wire [0:0] out_result_121__gfpga;
	wire [0:0] out_result_122__gfpga;
	wire [0:0] out_result_123__gfpga;
	wire [0:0] out_result_124__gfpga;
	wire [0:0] out_result_125__gfpga;
	wire [0:0] out_result_126__gfpga;
	wire [0:0] out_result_127__gfpga;

// ----- Benchmark outputs -------
	wire [0:0] out_result_0__bench;
	wire [0:0] out_result_1__bench;
	wire [0:0] out_result_2__bench;
	wire [0:0] out_result_3__bench;
	wire [0:0] out_result_4__bench;
	wire [0:0] out_result_5__bench;
	wire [0:0] out_result_6__bench;
	wire [0:0] out_result_7__bench;
	wire [0:0] out_result_8__bench;
	wire [0:0] out_result_9__bench;
	wire [0:0] out_result_10__bench;
	wire [0:0] out_result_11__bench;
	wire [0:0] out_result_12__bench;
	wire [0:0] out_result_13__bench;
	wire [0:0] out_result_14__bench;
	wire [0:0] out_result_15__bench;
	wire [0:0] out_result_16__bench;
	wire [0:0] out_result_17__bench;
	wire [0:0] out_result_18__bench;
	wire [0:0] out_result_19__bench;
	wire [0:0] out_result_20__bench;
	wire [0:0] out_result_21__bench;
	wire [0:0] out_result_22__bench;
	wire [0:0] out_result_23__bench;
	wire [0:0] out_result_24__bench;
	wire [0:0] out_result_25__bench;
	wire [0:0] out_result_26__bench;
	wire [0:0] out_result_27__bench;
	wire [0:0] out_result_28__bench;
	wire [0:0] out_result_29__bench;
	wire [0:0] out_result_30__bench;
	wire [0:0] out_result_31__bench;
	wire [0:0] out_result_32__bench;
	wire [0:0] out_result_33__bench;
	wire [0:0] out_result_34__bench;
	wire [0:0] out_result_35__bench;
	wire [0:0] out_result_36__bench;
	wire [0:0] out_result_37__bench;
	wire [0:0] out_result_38__bench;
	wire [0:0] out_result_39__bench;
	wire [0:0] out_result_40__bench;
	wire [0:0] out_result_41__bench;
	wire [0:0] out_result_42__bench;
	wire [0:0] out_result_43__bench;
	wire [0:0] out_result_44__bench;
	wire [0:0] out_result_45__bench;
	wire [0:0] out_result_46__bench;
	wire [0:0] out_result_47__bench;
	wire [0:0] out_result_48__bench;
	wire [0:0] out_result_49__bench;
	wire [0:0] out_result_50__bench;
	wire [0:0] out_result_51__bench;
	wire [0:0] out_result_52__bench;
	wire [0:0] out_result_53__bench;
	wire [0:0] out_result_54__bench;
	wire [0:0] out_result_55__bench;
	wire [0:0] out_result_56__bench;
	wire [0:0] out_result_57__bench;
	wire [0:0] out_result_58__bench;
	wire [0:0] out_result_59__bench;
	wire [0:0] out_result_60__bench;
	wire [0:0] out_result_61__bench;
	wire [0:0] out_result_62__bench;
	wire [0:0] out_result_63__bench;
	wire [0:0] out_result_64__bench;
	wire [0:0] out_result_65__bench;
	wire [0:0] out_result_66__bench;
	wire [0:0] out_result_67__bench;
	wire [0:0] out_result_68__bench;
	wire [0:0] out_result_69__bench;
	wire [0:0] out_result_70__bench;
	wire [0:0] out_result_71__bench;
	wire [0:0] out_result_72__bench;
	wire [0:0] out_result_73__bench;
	wire [0:0] out_result_74__bench;
	wire [0:0] out_result_75__bench;
	wire [0:0] out_result_76__bench;
	wire [0:0] out_result_77__bench;
	wire [0:0] out_result_78__bench;
	wire [0:0] out_result_79__bench;
	wire [0:0] out_result_80__bench;
	wire [0:0] out_result_81__bench;
	wire [0:0] out_result_82__bench;
	wire [0:0] out_result_83__bench;
	wire [0:0] out_result_84__bench;
	wire [0:0] out_result_85__bench;
	wire [0:0] out_result_86__bench;
	wire [0:0] out_result_87__bench;
	wire [0:0] out_result_88__bench;
	wire [0:0] out_result_89__bench;
	wire [0:0] out_result_90__bench;
	wire [0:0] out_result_91__bench;
	wire [0:0] out_result_92__bench;
	wire [0:0] out_result_93__bench;
	wire [0:0] out_result_94__bench;
	wire [0:0] out_result_95__bench;
	wire [0:0] out_result_96__bench;
	wire [0:0] out_result_97__bench;
	wire [0:0] out_result_98__bench;
	wire [0:0] out_result_99__bench;
	wire [0:0] out_result_100__bench;
	wire [0:0] out_result_101__bench;
	wire [0:0] out_result_102__bench;
	wire [0:0] out_result_103__bench;
	wire [0:0] out_result_104__bench;
	wire [0:0] out_result_105__bench;
	wire [0:0] out_result_106__bench;
	wire [0:0] out_result_107__bench;
	wire [0:0] out_result_108__bench;
	wire [0:0] out_result_109__bench;
	wire [0:0] out_result_110__bench;
	wire [0:0] out_result_111__bench;
	wire [0:0] out_result_112__bench;
	wire [0:0] out_result_113__bench;
	wire [0:0] out_result_114__bench;
	wire [0:0] out_result_115__bench;
	wire [0:0] out_result_116__bench;
	wire [0:0] out_result_117__bench;
	wire [0:0] out_result_118__bench;
	wire [0:0] out_result_119__bench;
	wire [0:0] out_result_120__bench;
	wire [0:0] out_result_121__bench;
	wire [0:0] out_result_122__bench;
	wire [0:0] out_result_123__bench;
	wire [0:0] out_result_124__bench;
	wire [0:0] out_result_125__bench;
	wire [0:0] out_result_126__bench;
	wire [0:0] out_result_127__bench;

// ----- Output vectors checking flags -------
	reg [0:0] out_result_0__flag;
	reg [0:0] out_result_1__flag;
	reg [0:0] out_result_2__flag;
	reg [0:0] out_result_3__flag;
	reg [0:0] out_result_4__flag;
	reg [0:0] out_result_5__flag;
	reg [0:0] out_result_6__flag;
	reg [0:0] out_result_7__flag;
	reg [0:0] out_result_8__flag;
	reg [0:0] out_result_9__flag;
	reg [0:0] out_result_10__flag;
	reg [0:0] out_result_11__flag;
	reg [0:0] out_result_12__flag;
	reg [0:0] out_result_13__flag;
	reg [0:0] out_result_14__flag;
	reg [0:0] out_result_15__flag;
	reg [0:0] out_result_16__flag;
	reg [0:0] out_result_17__flag;
	reg [0:0] out_result_18__flag;
	reg [0:0] out_result_19__flag;
	reg [0:0] out_result_20__flag;
	reg [0:0] out_result_21__flag;
	reg [0:0] out_result_22__flag;
	reg [0:0] out_result_23__flag;
	reg [0:0] out_result_24__flag;
	reg [0:0] out_result_25__flag;
	reg [0:0] out_result_26__flag;
	reg [0:0] out_result_27__flag;
	reg [0:0] out_result_28__flag;
	reg [0:0] out_result_29__flag;
	reg [0:0] out_result_30__flag;
	reg [0:0] out_result_31__flag;
	reg [0:0] out_result_32__flag;
	reg [0:0] out_result_33__flag;
	reg [0:0] out_result_34__flag;
	reg [0:0] out_result_35__flag;
	reg [0:0] out_result_36__flag;
	reg [0:0] out_result_37__flag;
	reg [0:0] out_result_38__flag;
	reg [0:0] out_result_39__flag;
	reg [0:0] out_result_40__flag;
	reg [0:0] out_result_41__flag;
	reg [0:0] out_result_42__flag;
	reg [0:0] out_result_43__flag;
	reg [0:0] out_result_44__flag;
	reg [0:0] out_result_45__flag;
	reg [0:0] out_result_46__flag;
	reg [0:0] out_result_47__flag;
	reg [0:0] out_result_48__flag;
	reg [0:0] out_result_49__flag;
	reg [0:0] out_result_50__flag;
	reg [0:0] out_result_51__flag;
	reg [0:0] out_result_52__flag;
	reg [0:0] out_result_53__flag;
	reg [0:0] out_result_54__flag;
	reg [0:0] out_result_55__flag;
	reg [0:0] out_result_56__flag;
	reg [0:0] out_result_57__flag;
	reg [0:0] out_result_58__flag;
	reg [0:0] out_result_59__flag;
	reg [0:0] out_result_60__flag;
	reg [0:0] out_result_61__flag;
	reg [0:0] out_result_62__flag;
	reg [0:0] out_result_63__flag;
	reg [0:0] out_result_64__flag;
	reg [0:0] out_result_65__flag;
	reg [0:0] out_result_66__flag;
	reg [0:0] out_result_67__flag;
	reg [0:0] out_result_68__flag;
	reg [0:0] out_result_69__flag;
	reg [0:0] out_result_70__flag;
	reg [0:0] out_result_71__flag;
	reg [0:0] out_result_72__flag;
	reg [0:0] out_result_73__flag;
	reg [0:0] out_result_74__flag;
	reg [0:0] out_result_75__flag;
	reg [0:0] out_result_76__flag;
	reg [0:0] out_result_77__flag;
	reg [0:0] out_result_78__flag;
	reg [0:0] out_result_79__flag;
	reg [0:0] out_result_80__flag;
	reg [0:0] out_result_81__flag;
	reg [0:0] out_result_82__flag;
	reg [0:0] out_result_83__flag;
	reg [0:0] out_result_84__flag;
	reg [0:0] out_result_85__flag;
	reg [0:0] out_result_86__flag;
	reg [0:0] out_result_87__flag;
	reg [0:0] out_result_88__flag;
	reg [0:0] out_result_89__flag;
	reg [0:0] out_result_90__flag;
	reg [0:0] out_result_91__flag;
	reg [0:0] out_result_92__flag;
	reg [0:0] out_result_93__flag;
	reg [0:0] out_result_94__flag;
	reg [0:0] out_result_95__flag;
	reg [0:0] out_result_96__flag;
	reg [0:0] out_result_97__flag;
	reg [0:0] out_result_98__flag;
	reg [0:0] out_result_99__flag;
	reg [0:0] out_result_100__flag;
	reg [0:0] out_result_101__flag;
	reg [0:0] out_result_102__flag;
	reg [0:0] out_result_103__flag;
	reg [0:0] out_result_104__flag;
	reg [0:0] out_result_105__flag;
	reg [0:0] out_result_106__flag;
	reg [0:0] out_result_107__flag;
	reg [0:0] out_result_108__flag;
	reg [0:0] out_result_109__flag;
	reg [0:0] out_result_110__flag;
	reg [0:0] out_result_111__flag;
	reg [0:0] out_result_112__flag;
	reg [0:0] out_result_113__flag;
	reg [0:0] out_result_114__flag;
	reg [0:0] out_result_115__flag;
	reg [0:0] out_result_116__flag;
	reg [0:0] out_result_117__flag;
	reg [0:0] out_result_118__flag;
	reg [0:0] out_result_119__flag;
	reg [0:0] out_result_120__flag;
	reg [0:0] out_result_121__flag;
	reg [0:0] out_result_122__flag;
	reg [0:0] out_result_123__flag;
	reg [0:0] out_result_124__flag;
	reg [0:0] out_result_125__flag;
	reg [0:0] out_result_126__flag;
	reg [0:0] out_result_127__flag;

// ----- Error counter -------
	integer nb_error= 0;

// ----- FPGA fabric instanciation -------
	counter_top_formal_verification FPGA_DUT(
		clk,
		resetb,
		out_result_0__gfpga,
		out_result_1__gfpga,
		out_result_2__gfpga,
		out_result_3__gfpga,
		out_result_4__gfpga,
		out_result_5__gfpga,
		out_result_6__gfpga,
		out_result_7__gfpga,
		out_result_8__gfpga,
		out_result_9__gfpga,
		out_result_10__gfpga,
		out_result_11__gfpga,
		out_result_12__gfpga,
		out_result_13__gfpga,
		out_result_14__gfpga,
		out_result_15__gfpga,
		out_result_16__gfpga,
		out_result_17__gfpga,
		out_result_18__gfpga,
		out_result_19__gfpga,
		out_result_20__gfpga,
		out_result_21__gfpga,
		out_result_22__gfpga,
		out_result_23__gfpga,
		out_result_24__gfpga,
		out_result_25__gfpga,
		out_result_26__gfpga,
		out_result_27__gfpga,
		out_result_28__gfpga,
		out_result_29__gfpga,
		out_result_30__gfpga,
		out_result_31__gfpga,
		out_result_32__gfpga,
		out_result_33__gfpga,
		out_result_34__gfpga,
		out_result_35__gfpga,
		out_result_36__gfpga,
		out_result_37__gfpga,
		out_result_38__gfpga,
		out_result_39__gfpga,
		out_result_40__gfpga,
		out_result_41__gfpga,
		out_result_42__gfpga,
		out_result_43__gfpga,
		out_result_44__gfpga,
		out_result_45__gfpga,
		out_result_46__gfpga,
		out_result_47__gfpga,
		out_result_48__gfpga,
		out_result_49__gfpga,
		out_result_50__gfpga,
		out_result_51__gfpga,
		out_result_52__gfpga,
		out_result_53__gfpga,
		out_result_54__gfpga,
		out_result_55__gfpga,
		out_result_56__gfpga,
		out_result_57__gfpga,
		out_result_58__gfpga,
		out_result_59__gfpga,
		out_result_60__gfpga,
		out_result_61__gfpga,
		out_result_62__gfpga,
		out_result_63__gfpga,
		out_result_64__gfpga,
		out_result_65__gfpga,
		out_result_66__gfpga,
		out_result_67__gfpga,
		out_result_68__gfpga,
		out_result_69__gfpga,
		out_result_70__gfpga,
		out_result_71__gfpga,
		out_result_72__gfpga,
		out_result_73__gfpga,
		out_result_74__gfpga,
		out_result_75__gfpga,
		out_result_76__gfpga,
		out_result_77__gfpga,
		out_result_78__gfpga,
		out_result_79__gfpga,
		out_result_80__gfpga,
		out_result_81__gfpga,
		out_result_82__gfpga,
		out_result_83__gfpga,
		out_result_84__gfpga,
		out_result_85__gfpga,
		out_result_86__gfpga,
		out_result_87__gfpga,
		out_result_88__gfpga,
		out_result_89__gfpga,
		out_result_90__gfpga,
		out_result_91__gfpga,
		out_result_92__gfpga,
		out_result_93__gfpga,
		out_result_94__gfpga,
		out_result_95__gfpga,
		out_result_96__gfpga,
		out_result_97__gfpga,
		out_result_98__gfpga,
		out_result_99__gfpga,
		out_result_100__gfpga,
		out_result_101__gfpga,
		out_result_102__gfpga,
		out_result_103__gfpga,
		out_result_104__gfpga,
		out_result_105__gfpga,
		out_result_106__gfpga,
		out_result_107__gfpga,
		out_result_108__gfpga,
		out_result_109__gfpga,
		out_result_110__gfpga,
		out_result_111__gfpga,
		out_result_112__gfpga,
		out_result_113__gfpga,
		out_result_114__gfpga,
		out_result_115__gfpga,
		out_result_116__gfpga,
		out_result_117__gfpga,
		out_result_118__gfpga,
		out_result_119__gfpga,
		out_result_120__gfpga,
		out_result_121__gfpga,
		out_result_122__gfpga,
		out_result_123__gfpga,
		out_result_124__gfpga,
		out_result_125__gfpga,
		out_result_126__gfpga,
		out_result_127__gfpga	);
// ----- End FPGA Fabric Instanication -------

// ----- Reference Benchmark Instanication -------
	counter REF_DUT(
		clk,
		resetb,
		out_result_0__bench,
		out_result_1__bench,
		out_result_2__bench,
		out_result_3__bench,
		out_result_4__bench,
		out_result_5__bench,
		out_result_6__bench,
		out_result_7__bench,
		out_result_8__bench,
		out_result_9__bench,
		out_result_10__bench,
		out_result_11__bench,
		out_result_12__bench,
		out_result_13__bench,
		out_result_14__bench,
		out_result_15__bench,
		out_result_16__bench,
		out_result_17__bench,
		out_result_18__bench,
		out_result_19__bench,
		out_result_20__bench,
		out_result_21__bench,
		out_result_22__bench,
		out_result_23__bench,
		out_result_24__bench,
		out_result_25__bench,
		out_result_26__bench,
		out_result_27__bench,
		out_result_28__bench,
		out_result_29__bench,
		out_result_30__bench,
		out_result_31__bench,
		out_result_32__bench,
		out_result_33__bench,
		out_result_34__bench,
		out_result_35__bench,
		out_result_36__bench,
		out_result_37__bench,
		out_result_38__bench,
		out_result_39__bench,
		out_result_40__bench,
		out_result_41__bench,
		out_result_42__bench,
		out_result_43__bench,
		out_result_44__bench,
		out_result_45__bench,
		out_result_46__bench,
		out_result_47__bench,
		out_result_48__bench,
		out_result_49__bench,
		out_result_50__bench,
		out_result_51__bench,
		out_result_52__bench,
		out_result_53__bench,
		out_result_54__bench,
		out_result_55__bench,
		out_result_56__bench,
		out_result_57__bench,
		out_result_58__bench,
		out_result_59__bench,
		out_result_60__bench,
		out_result_61__bench,
		out_result_62__bench,
		out_result_63__bench,
		out_result_64__bench,
		out_result_65__bench,
		out_result_66__bench,
		out_result_67__bench,
		out_result_68__bench,
		out_result_69__bench,
		out_result_70__bench,
		out_result_71__bench,
		out_result_72__bench,
		out_result_73__bench,
		out_result_74__bench,
		out_result_75__bench,
		out_result_76__bench,
		out_result_77__bench,
		out_result_78__bench,
		out_result_79__bench,
		out_result_80__bench,
		out_result_81__bench,
		out_result_82__bench,
		out_result_83__bench,
		out_result_84__bench,
		out_result_85__bench,
		out_result_86__bench,
		out_result_87__bench,
		out_result_88__bench,
		out_result_89__bench,
		out_result_90__bench,
		out_result_91__bench,
		out_result_92__bench,
		out_result_93__bench,
		out_result_94__bench,
		out_result_95__bench,
		out_result_96__bench,
		out_result_97__bench,
		out_result_98__bench,
		out_result_99__bench,
		out_result_100__bench,
		out_result_101__bench,
		out_result_102__bench,
		out_result_103__bench,
		out_result_104__bench,
		out_result_105__bench,
		out_result_106__bench,
		out_result_107__bench,
		out_result_108__bench,
		out_result_109__bench,
		out_result_110__bench,
		out_result_111__bench,
		out_result_112__bench,
		out_result_113__bench,
		out_result_114__bench,
		out_result_115__bench,
		out_result_116__bench,
		out_result_117__bench,
		out_result_118__bench,
		out_result_119__bench,
		out_result_120__bench,
		out_result_121__bench,
		out_result_122__bench,
		out_result_123__bench,
		out_result_124__bench,
		out_result_125__bench,
		out_result_126__bench,
		out_result_127__bench	);
// ----- End reference Benchmark Instanication -------

// ----- Clock 'clk' Initialization -------
	initial begin
		clk[0] <= 1'b0;
		while(1) begin
			#1
			clk[0] <= !clk[0];
		end
	end

// ----- Begin reset signal generation -----
// ----- End reset signal generation -----

// ----- Input Initialization -------
	initial begin
		resetb <= 1'b0;

		out_result_0__flag[0] <= 1'b0;
		out_result_1__flag[0] <= 1'b0;
		out_result_2__flag[0] <= 1'b0;
		out_result_3__flag[0] <= 1'b0;
		out_result_4__flag[0] <= 1'b0;
		out_result_5__flag[0] <= 1'b0;
		out_result_6__flag[0] <= 1'b0;
		out_result_7__flag[0] <= 1'b0;
		out_result_8__flag[0] <= 1'b0;
		out_result_9__flag[0] <= 1'b0;
		out_result_10__flag[0] <= 1'b0;
		out_result_11__flag[0] <= 1'b0;
		out_result_12__flag[0] <= 1'b0;
		out_result_13__flag[0] <= 1'b0;
		out_result_14__flag[0] <= 1'b0;
		out_result_15__flag[0] <= 1'b0;
		out_result_16__flag[0] <= 1'b0;
		out_result_17__flag[0] <= 1'b0;
		out_result_18__flag[0] <= 1'b0;
		out_result_19__flag[0] <= 1'b0;
		out_result_20__flag[0] <= 1'b0;
		out_result_21__flag[0] <= 1'b0;
		out_result_22__flag[0] <= 1'b0;
		out_result_23__flag[0] <= 1'b0;
		out_result_24__flag[0] <= 1'b0;
		out_result_25__flag[0] <= 1'b0;
		out_result_26__flag[0] <= 1'b0;
		out_result_27__flag[0] <= 1'b0;
		out_result_28__flag[0] <= 1'b0;
		out_result_29__flag[0] <= 1'b0;
		out_result_30__flag[0] <= 1'b0;
		out_result_31__flag[0] <= 1'b0;
		out_result_32__flag[0] <= 1'b0;
		out_result_33__flag[0] <= 1'b0;
		out_result_34__flag[0] <= 1'b0;
		out_result_35__flag[0] <= 1'b0;
		out_result_36__flag[0] <= 1'b0;
		out_result_37__flag[0] <= 1'b0;
		out_result_38__flag[0] <= 1'b0;
		out_result_39__flag[0] <= 1'b0;
		out_result_40__flag[0] <= 1'b0;
		out_result_41__flag[0] <= 1'b0;
		out_result_42__flag[0] <= 1'b0;
		out_result_43__flag[0] <= 1'b0;
		out_result_44__flag[0] <= 1'b0;
		out_result_45__flag[0] <= 1'b0;
		out_result_46__flag[0] <= 1'b0;
		out_result_47__flag[0] <= 1'b0;
		out_result_48__flag[0] <= 1'b0;
		out_result_49__flag[0] <= 1'b0;
		out_result_50__flag[0] <= 1'b0;
		out_result_51__flag[0] <= 1'b0;
		out_result_52__flag[0] <= 1'b0;
		out_result_53__flag[0] <= 1'b0;
		out_result_54__flag[0] <= 1'b0;
		out_result_55__flag[0] <= 1'b0;
		out_result_56__flag[0] <= 1'b0;
		out_result_57__flag[0] <= 1'b0;
		out_result_58__flag[0] <= 1'b0;
		out_result_59__flag[0] <= 1'b0;
		out_result_60__flag[0] <= 1'b0;
		out_result_61__flag[0] <= 1'b0;
		out_result_62__flag[0] <= 1'b0;
		out_result_63__flag[0] <= 1'b0;
		out_result_64__flag[0] <= 1'b0;
		out_result_65__flag[0] <= 1'b0;
		out_result_66__flag[0] <= 1'b0;
		out_result_67__flag[0] <= 1'b0;
		out_result_68__flag[0] <= 1'b0;
		out_result_69__flag[0] <= 1'b0;
		out_result_70__flag[0] <= 1'b0;
		out_result_71__flag[0] <= 1'b0;
		out_result_72__flag[0] <= 1'b0;
		out_result_73__flag[0] <= 1'b0;
		out_result_74__flag[0] <= 1'b0;
		out_result_75__flag[0] <= 1'b0;
		out_result_76__flag[0] <= 1'b0;
		out_result_77__flag[0] <= 1'b0;
		out_result_78__flag[0] <= 1'b0;
		out_result_79__flag[0] <= 1'b0;
		out_result_80__flag[0] <= 1'b0;
		out_result_81__flag[0] <= 1'b0;
		out_result_82__flag[0] <= 1'b0;
		out_result_83__flag[0] <= 1'b0;
		out_result_84__flag[0] <= 1'b0;
		out_result_85__flag[0] <= 1'b0;
		out_result_86__flag[0] <= 1'b0;
		out_result_87__flag[0] <= 1'b0;
		out_result_88__flag[0] <= 1'b0;
		out_result_89__flag[0] <= 1'b0;
		out_result_90__flag[0] <= 1'b0;
		out_result_91__flag[0] <= 1'b0;
		out_result_92__flag[0] <= 1'b0;
		out_result_93__flag[0] <= 1'b0;
		out_result_94__flag[0] <= 1'b0;
		out_result_95__flag[0] <= 1'b0;
		out_result_96__flag[0] <= 1'b0;
		out_result_97__flag[0] <= 1'b0;
		out_result_98__flag[0] <= 1'b0;
		out_result_99__flag[0] <= 1'b0;
		out_result_100__flag[0] <= 1'b0;
		out_result_101__flag[0] <= 1'b0;
		out_result_102__flag[0] <= 1'b0;
		out_result_103__flag[0] <= 1'b0;
		out_result_104__flag[0] <= 1'b0;
		out_result_105__flag[0] <= 1'b0;
		out_result_106__flag[0] <= 1'b0;
		out_result_107__flag[0] <= 1'b0;
		out_result_108__flag[0] <= 1'b0;
		out_result_109__flag[0] <= 1'b0;
		out_result_110__flag[0] <= 1'b0;
		out_result_111__flag[0] <= 1'b0;
		out_result_112__flag[0] <= 1'b0;
		out_result_113__flag[0] <= 1'b0;
		out_result_114__flag[0] <= 1'b0;
		out_result_115__flag[0] <= 1'b0;
		out_result_116__flag[0] <= 1'b0;
		out_result_117__flag[0] <= 1'b0;
		out_result_118__flag[0] <= 1'b0;
		out_result_119__flag[0] <= 1'b0;
		out_result_120__flag[0] <= 1'b0;
		out_result_121__flag[0] <= 1'b0;
		out_result_122__flag[0] <= 1'b0;
		out_result_123__flag[0] <= 1'b0;
		out_result_124__flag[0] <= 1'b0;
		out_result_125__flag[0] <= 1'b0;
		out_result_126__flag[0] <= 1'b0;
		out_result_127__flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge clk[0]) begin
		resetb <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge clk[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else begin
			if(!(out_result_0__gfpga === out_result_0__bench) && !(out_result_0__bench === 1'bx)) begin
				out_result_0__flag <= 1'b1;
			end else begin
				out_result_0__flag<= 1'b0;
			end
			if(!(out_result_1__gfpga === out_result_1__bench) && !(out_result_1__bench === 1'bx)) begin
				out_result_1__flag <= 1'b1;
			end else begin
				out_result_1__flag<= 1'b0;
			end
			if(!(out_result_2__gfpga === out_result_2__bench) && !(out_result_2__bench === 1'bx)) begin
				out_result_2__flag <= 1'b1;
			end else begin
				out_result_2__flag<= 1'b0;
			end
			if(!(out_result_3__gfpga === out_result_3__bench) && !(out_result_3__bench === 1'bx)) begin
				out_result_3__flag <= 1'b1;
			end else begin
				out_result_3__flag<= 1'b0;
			end
			if(!(out_result_4__gfpga === out_result_4__bench) && !(out_result_4__bench === 1'bx)) begin
				out_result_4__flag <= 1'b1;
			end else begin
				out_result_4__flag<= 1'b0;
			end
			if(!(out_result_5__gfpga === out_result_5__bench) && !(out_result_5__bench === 1'bx)) begin
				out_result_5__flag <= 1'b1;
			end else begin
				out_result_5__flag<= 1'b0;
			end
			if(!(out_result_6__gfpga === out_result_6__bench) && !(out_result_6__bench === 1'bx)) begin
				out_result_6__flag <= 1'b1;
			end else begin
				out_result_6__flag<= 1'b0;
			end
			if(!(out_result_7__gfpga === out_result_7__bench) && !(out_result_7__bench === 1'bx)) begin
				out_result_7__flag <= 1'b1;
			end else begin
				out_result_7__flag<= 1'b0;
			end
			if(!(out_result_8__gfpga === out_result_8__bench) && !(out_result_8__bench === 1'bx)) begin
				out_result_8__flag <= 1'b1;
			end else begin
				out_result_8__flag<= 1'b0;
			end
			if(!(out_result_9__gfpga === out_result_9__bench) && !(out_result_9__bench === 1'bx)) begin
				out_result_9__flag <= 1'b1;
			end else begin
				out_result_9__flag<= 1'b0;
			end
			if(!(out_result_10__gfpga === out_result_10__bench) && !(out_result_10__bench === 1'bx)) begin
				out_result_10__flag <= 1'b1;
			end else begin
				out_result_10__flag<= 1'b0;
			end
			if(!(out_result_11__gfpga === out_result_11__bench) && !(out_result_11__bench === 1'bx)) begin
				out_result_11__flag <= 1'b1;
			end else begin
				out_result_11__flag<= 1'b0;
			end
			if(!(out_result_12__gfpga === out_result_12__bench) && !(out_result_12__bench === 1'bx)) begin
				out_result_12__flag <= 1'b1;
			end else begin
				out_result_12__flag<= 1'b0;
			end
			if(!(out_result_13__gfpga === out_result_13__bench) && !(out_result_13__bench === 1'bx)) begin
				out_result_13__flag <= 1'b1;
			end else begin
				out_result_13__flag<= 1'b0;
			end
			if(!(out_result_14__gfpga === out_result_14__bench) && !(out_result_14__bench === 1'bx)) begin
				out_result_14__flag <= 1'b1;
			end else begin
				out_result_14__flag<= 1'b0;
			end
			if(!(out_result_15__gfpga === out_result_15__bench) && !(out_result_15__bench === 1'bx)) begin
				out_result_15__flag <= 1'b1;
			end else begin
				out_result_15__flag<= 1'b0;
			end
			if(!(out_result_16__gfpga === out_result_16__bench) && !(out_result_16__bench === 1'bx)) begin
				out_result_16__flag <= 1'b1;
			end else begin
				out_result_16__flag<= 1'b0;
			end
			if(!(out_result_17__gfpga === out_result_17__bench) && !(out_result_17__bench === 1'bx)) begin
				out_result_17__flag <= 1'b1;
			end else begin
				out_result_17__flag<= 1'b0;
			end
			if(!(out_result_18__gfpga === out_result_18__bench) && !(out_result_18__bench === 1'bx)) begin
				out_result_18__flag <= 1'b1;
			end else begin
				out_result_18__flag<= 1'b0;
			end
			if(!(out_result_19__gfpga === out_result_19__bench) && !(out_result_19__bench === 1'bx)) begin
				out_result_19__flag <= 1'b1;
			end else begin
				out_result_19__flag<= 1'b0;
			end
			if(!(out_result_20__gfpga === out_result_20__bench) && !(out_result_20__bench === 1'bx)) begin
				out_result_20__flag <= 1'b1;
			end else begin
				out_result_20__flag<= 1'b0;
			end
			if(!(out_result_21__gfpga === out_result_21__bench) && !(out_result_21__bench === 1'bx)) begin
				out_result_21__flag <= 1'b1;
			end else begin
				out_result_21__flag<= 1'b0;
			end
			if(!(out_result_22__gfpga === out_result_22__bench) && !(out_result_22__bench === 1'bx)) begin
				out_result_22__flag <= 1'b1;
			end else begin
				out_result_22__flag<= 1'b0;
			end
			if(!(out_result_23__gfpga === out_result_23__bench) && !(out_result_23__bench === 1'bx)) begin
				out_result_23__flag <= 1'b1;
			end else begin
				out_result_23__flag<= 1'b0;
			end
			if(!(out_result_24__gfpga === out_result_24__bench) && !(out_result_24__bench === 1'bx)) begin
				out_result_24__flag <= 1'b1;
			end else begin
				out_result_24__flag<= 1'b0;
			end
			if(!(out_result_25__gfpga === out_result_25__bench) && !(out_result_25__bench === 1'bx)) begin
				out_result_25__flag <= 1'b1;
			end else begin
				out_result_25__flag<= 1'b0;
			end
			if(!(out_result_26__gfpga === out_result_26__bench) && !(out_result_26__bench === 1'bx)) begin
				out_result_26__flag <= 1'b1;
			end else begin
				out_result_26__flag<= 1'b0;
			end
			if(!(out_result_27__gfpga === out_result_27__bench) && !(out_result_27__bench === 1'bx)) begin
				out_result_27__flag <= 1'b1;
			end else begin
				out_result_27__flag<= 1'b0;
			end
			if(!(out_result_28__gfpga === out_result_28__bench) && !(out_result_28__bench === 1'bx)) begin
				out_result_28__flag <= 1'b1;
			end else begin
				out_result_28__flag<= 1'b0;
			end
			if(!(out_result_29__gfpga === out_result_29__bench) && !(out_result_29__bench === 1'bx)) begin
				out_result_29__flag <= 1'b1;
			end else begin
				out_result_29__flag<= 1'b0;
			end
			if(!(out_result_30__gfpga === out_result_30__bench) && !(out_result_30__bench === 1'bx)) begin
				out_result_30__flag <= 1'b1;
			end else begin
				out_result_30__flag<= 1'b0;
			end
			if(!(out_result_31__gfpga === out_result_31__bench) && !(out_result_31__bench === 1'bx)) begin
				out_result_31__flag <= 1'b1;
			end else begin
				out_result_31__flag<= 1'b0;
			end
			if(!(out_result_32__gfpga === out_result_32__bench) && !(out_result_32__bench === 1'bx)) begin
				out_result_32__flag <= 1'b1;
			end else begin
				out_result_32__flag<= 1'b0;
			end
			if(!(out_result_33__gfpga === out_result_33__bench) && !(out_result_33__bench === 1'bx)) begin
				out_result_33__flag <= 1'b1;
			end else begin
				out_result_33__flag<= 1'b0;
			end
			if(!(out_result_34__gfpga === out_result_34__bench) && !(out_result_34__bench === 1'bx)) begin
				out_result_34__flag <= 1'b1;
			end else begin
				out_result_34__flag<= 1'b0;
			end
			if(!(out_result_35__gfpga === out_result_35__bench) && !(out_result_35__bench === 1'bx)) begin
				out_result_35__flag <= 1'b1;
			end else begin
				out_result_35__flag<= 1'b0;
			end
			if(!(out_result_36__gfpga === out_result_36__bench) && !(out_result_36__bench === 1'bx)) begin
				out_result_36__flag <= 1'b1;
			end else begin
				out_result_36__flag<= 1'b0;
			end
			if(!(out_result_37__gfpga === out_result_37__bench) && !(out_result_37__bench === 1'bx)) begin
				out_result_37__flag <= 1'b1;
			end else begin
				out_result_37__flag<= 1'b0;
			end
			if(!(out_result_38__gfpga === out_result_38__bench) && !(out_result_38__bench === 1'bx)) begin
				out_result_38__flag <= 1'b1;
			end else begin
				out_result_38__flag<= 1'b0;
			end
			if(!(out_result_39__gfpga === out_result_39__bench) && !(out_result_39__bench === 1'bx)) begin
				out_result_39__flag <= 1'b1;
			end else begin
				out_result_39__flag<= 1'b0;
			end
			if(!(out_result_40__gfpga === out_result_40__bench) && !(out_result_40__bench === 1'bx)) begin
				out_result_40__flag <= 1'b1;
			end else begin
				out_result_40__flag<= 1'b0;
			end
			if(!(out_result_41__gfpga === out_result_41__bench) && !(out_result_41__bench === 1'bx)) begin
				out_result_41__flag <= 1'b1;
			end else begin
				out_result_41__flag<= 1'b0;
			end
			if(!(out_result_42__gfpga === out_result_42__bench) && !(out_result_42__bench === 1'bx)) begin
				out_result_42__flag <= 1'b1;
			end else begin
				out_result_42__flag<= 1'b0;
			end
			if(!(out_result_43__gfpga === out_result_43__bench) && !(out_result_43__bench === 1'bx)) begin
				out_result_43__flag <= 1'b1;
			end else begin
				out_result_43__flag<= 1'b0;
			end
			if(!(out_result_44__gfpga === out_result_44__bench) && !(out_result_44__bench === 1'bx)) begin
				out_result_44__flag <= 1'b1;
			end else begin
				out_result_44__flag<= 1'b0;
			end
			if(!(out_result_45__gfpga === out_result_45__bench) && !(out_result_45__bench === 1'bx)) begin
				out_result_45__flag <= 1'b1;
			end else begin
				out_result_45__flag<= 1'b0;
			end
			if(!(out_result_46__gfpga === out_result_46__bench) && !(out_result_46__bench === 1'bx)) begin
				out_result_46__flag <= 1'b1;
			end else begin
				out_result_46__flag<= 1'b0;
			end
			if(!(out_result_47__gfpga === out_result_47__bench) && !(out_result_47__bench === 1'bx)) begin
				out_result_47__flag <= 1'b1;
			end else begin
				out_result_47__flag<= 1'b0;
			end
			if(!(out_result_48__gfpga === out_result_48__bench) && !(out_result_48__bench === 1'bx)) begin
				out_result_48__flag <= 1'b1;
			end else begin
				out_result_48__flag<= 1'b0;
			end
			if(!(out_result_49__gfpga === out_result_49__bench) && !(out_result_49__bench === 1'bx)) begin
				out_result_49__flag <= 1'b1;
			end else begin
				out_result_49__flag<= 1'b0;
			end
			if(!(out_result_50__gfpga === out_result_50__bench) && !(out_result_50__bench === 1'bx)) begin
				out_result_50__flag <= 1'b1;
			end else begin
				out_result_50__flag<= 1'b0;
			end
			if(!(out_result_51__gfpga === out_result_51__bench) && !(out_result_51__bench === 1'bx)) begin
				out_result_51__flag <= 1'b1;
			end else begin
				out_result_51__flag<= 1'b0;
			end
			if(!(out_result_52__gfpga === out_result_52__bench) && !(out_result_52__bench === 1'bx)) begin
				out_result_52__flag <= 1'b1;
			end else begin
				out_result_52__flag<= 1'b0;
			end
			if(!(out_result_53__gfpga === out_result_53__bench) && !(out_result_53__bench === 1'bx)) begin
				out_result_53__flag <= 1'b1;
			end else begin
				out_result_53__flag<= 1'b0;
			end
			if(!(out_result_54__gfpga === out_result_54__bench) && !(out_result_54__bench === 1'bx)) begin
				out_result_54__flag <= 1'b1;
			end else begin
				out_result_54__flag<= 1'b0;
			end
			if(!(out_result_55__gfpga === out_result_55__bench) && !(out_result_55__bench === 1'bx)) begin
				out_result_55__flag <= 1'b1;
			end else begin
				out_result_55__flag<= 1'b0;
			end
			if(!(out_result_56__gfpga === out_result_56__bench) && !(out_result_56__bench === 1'bx)) begin
				out_result_56__flag <= 1'b1;
			end else begin
				out_result_56__flag<= 1'b0;
			end
			if(!(out_result_57__gfpga === out_result_57__bench) && !(out_result_57__bench === 1'bx)) begin
				out_result_57__flag <= 1'b1;
			end else begin
				out_result_57__flag<= 1'b0;
			end
			if(!(out_result_58__gfpga === out_result_58__bench) && !(out_result_58__bench === 1'bx)) begin
				out_result_58__flag <= 1'b1;
			end else begin
				out_result_58__flag<= 1'b0;
			end
			if(!(out_result_59__gfpga === out_result_59__bench) && !(out_result_59__bench === 1'bx)) begin
				out_result_59__flag <= 1'b1;
			end else begin
				out_result_59__flag<= 1'b0;
			end
			if(!(out_result_60__gfpga === out_result_60__bench) && !(out_result_60__bench === 1'bx)) begin
				out_result_60__flag <= 1'b1;
			end else begin
				out_result_60__flag<= 1'b0;
			end
			if(!(out_result_61__gfpga === out_result_61__bench) && !(out_result_61__bench === 1'bx)) begin
				out_result_61__flag <= 1'b1;
			end else begin
				out_result_61__flag<= 1'b0;
			end
			if(!(out_result_62__gfpga === out_result_62__bench) && !(out_result_62__bench === 1'bx)) begin
				out_result_62__flag <= 1'b1;
			end else begin
				out_result_62__flag<= 1'b0;
			end
			if(!(out_result_63__gfpga === out_result_63__bench) && !(out_result_63__bench === 1'bx)) begin
				out_result_63__flag <= 1'b1;
			end else begin
				out_result_63__flag<= 1'b0;
			end
			if(!(out_result_64__gfpga === out_result_64__bench) && !(out_result_64__bench === 1'bx)) begin
				out_result_64__flag <= 1'b1;
			end else begin
				out_result_64__flag<= 1'b0;
			end
			if(!(out_result_65__gfpga === out_result_65__bench) && !(out_result_65__bench === 1'bx)) begin
				out_result_65__flag <= 1'b1;
			end else begin
				out_result_65__flag<= 1'b0;
			end
			if(!(out_result_66__gfpga === out_result_66__bench) && !(out_result_66__bench === 1'bx)) begin
				out_result_66__flag <= 1'b1;
			end else begin
				out_result_66__flag<= 1'b0;
			end
			if(!(out_result_67__gfpga === out_result_67__bench) && !(out_result_67__bench === 1'bx)) begin
				out_result_67__flag <= 1'b1;
			end else begin
				out_result_67__flag<= 1'b0;
			end
			if(!(out_result_68__gfpga === out_result_68__bench) && !(out_result_68__bench === 1'bx)) begin
				out_result_68__flag <= 1'b1;
			end else begin
				out_result_68__flag<= 1'b0;
			end
			if(!(out_result_69__gfpga === out_result_69__bench) && !(out_result_69__bench === 1'bx)) begin
				out_result_69__flag <= 1'b1;
			end else begin
				out_result_69__flag<= 1'b0;
			end
			if(!(out_result_70__gfpga === out_result_70__bench) && !(out_result_70__bench === 1'bx)) begin
				out_result_70__flag <= 1'b1;
			end else begin
				out_result_70__flag<= 1'b0;
			end
			if(!(out_result_71__gfpga === out_result_71__bench) && !(out_result_71__bench === 1'bx)) begin
				out_result_71__flag <= 1'b1;
			end else begin
				out_result_71__flag<= 1'b0;
			end
			if(!(out_result_72__gfpga === out_result_72__bench) && !(out_result_72__bench === 1'bx)) begin
				out_result_72__flag <= 1'b1;
			end else begin
				out_result_72__flag<= 1'b0;
			end
			if(!(out_result_73__gfpga === out_result_73__bench) && !(out_result_73__bench === 1'bx)) begin
				out_result_73__flag <= 1'b1;
			end else begin
				out_result_73__flag<= 1'b0;
			end
			if(!(out_result_74__gfpga === out_result_74__bench) && !(out_result_74__bench === 1'bx)) begin
				out_result_74__flag <= 1'b1;
			end else begin
				out_result_74__flag<= 1'b0;
			end
			if(!(out_result_75__gfpga === out_result_75__bench) && !(out_result_75__bench === 1'bx)) begin
				out_result_75__flag <= 1'b1;
			end else begin
				out_result_75__flag<= 1'b0;
			end
			if(!(out_result_76__gfpga === out_result_76__bench) && !(out_result_76__bench === 1'bx)) begin
				out_result_76__flag <= 1'b1;
			end else begin
				out_result_76__flag<= 1'b0;
			end
			if(!(out_result_77__gfpga === out_result_77__bench) && !(out_result_77__bench === 1'bx)) begin
				out_result_77__flag <= 1'b1;
			end else begin
				out_result_77__flag<= 1'b0;
			end
			if(!(out_result_78__gfpga === out_result_78__bench) && !(out_result_78__bench === 1'bx)) begin
				out_result_78__flag <= 1'b1;
			end else begin
				out_result_78__flag<= 1'b0;
			end
			if(!(out_result_79__gfpga === out_result_79__bench) && !(out_result_79__bench === 1'bx)) begin
				out_result_79__flag <= 1'b1;
			end else begin
				out_result_79__flag<= 1'b0;
			end
			if(!(out_result_80__gfpga === out_result_80__bench) && !(out_result_80__bench === 1'bx)) begin
				out_result_80__flag <= 1'b1;
			end else begin
				out_result_80__flag<= 1'b0;
			end
			if(!(out_result_81__gfpga === out_result_81__bench) && !(out_result_81__bench === 1'bx)) begin
				out_result_81__flag <= 1'b1;
			end else begin
				out_result_81__flag<= 1'b0;
			end
			if(!(out_result_82__gfpga === out_result_82__bench) && !(out_result_82__bench === 1'bx)) begin
				out_result_82__flag <= 1'b1;
			end else begin
				out_result_82__flag<= 1'b0;
			end
			if(!(out_result_83__gfpga === out_result_83__bench) && !(out_result_83__bench === 1'bx)) begin
				out_result_83__flag <= 1'b1;
			end else begin
				out_result_83__flag<= 1'b0;
			end
			if(!(out_result_84__gfpga === out_result_84__bench) && !(out_result_84__bench === 1'bx)) begin
				out_result_84__flag <= 1'b1;
			end else begin
				out_result_84__flag<= 1'b0;
			end
			if(!(out_result_85__gfpga === out_result_85__bench) && !(out_result_85__bench === 1'bx)) begin
				out_result_85__flag <= 1'b1;
			end else begin
				out_result_85__flag<= 1'b0;
			end
			if(!(out_result_86__gfpga === out_result_86__bench) && !(out_result_86__bench === 1'bx)) begin
				out_result_86__flag <= 1'b1;
			end else begin
				out_result_86__flag<= 1'b0;
			end
			if(!(out_result_87__gfpga === out_result_87__bench) && !(out_result_87__bench === 1'bx)) begin
				out_result_87__flag <= 1'b1;
			end else begin
				out_result_87__flag<= 1'b0;
			end
			if(!(out_result_88__gfpga === out_result_88__bench) && !(out_result_88__bench === 1'bx)) begin
				out_result_88__flag <= 1'b1;
			end else begin
				out_result_88__flag<= 1'b0;
			end
			if(!(out_result_89__gfpga === out_result_89__bench) && !(out_result_89__bench === 1'bx)) begin
				out_result_89__flag <= 1'b1;
			end else begin
				out_result_89__flag<= 1'b0;
			end
			if(!(out_result_90__gfpga === out_result_90__bench) && !(out_result_90__bench === 1'bx)) begin
				out_result_90__flag <= 1'b1;
			end else begin
				out_result_90__flag<= 1'b0;
			end
			if(!(out_result_91__gfpga === out_result_91__bench) && !(out_result_91__bench === 1'bx)) begin
				out_result_91__flag <= 1'b1;
			end else begin
				out_result_91__flag<= 1'b0;
			end
			if(!(out_result_92__gfpga === out_result_92__bench) && !(out_result_92__bench === 1'bx)) begin
				out_result_92__flag <= 1'b1;
			end else begin
				out_result_92__flag<= 1'b0;
			end
			if(!(out_result_93__gfpga === out_result_93__bench) && !(out_result_93__bench === 1'bx)) begin
				out_result_93__flag <= 1'b1;
			end else begin
				out_result_93__flag<= 1'b0;
			end
			if(!(out_result_94__gfpga === out_result_94__bench) && !(out_result_94__bench === 1'bx)) begin
				out_result_94__flag <= 1'b1;
			end else begin
				out_result_94__flag<= 1'b0;
			end
			if(!(out_result_95__gfpga === out_result_95__bench) && !(out_result_95__bench === 1'bx)) begin
				out_result_95__flag <= 1'b1;
			end else begin
				out_result_95__flag<= 1'b0;
			end
			if(!(out_result_96__gfpga === out_result_96__bench) && !(out_result_96__bench === 1'bx)) begin
				out_result_96__flag <= 1'b1;
			end else begin
				out_result_96__flag<= 1'b0;
			end
			if(!(out_result_97__gfpga === out_result_97__bench) && !(out_result_97__bench === 1'bx)) begin
				out_result_97__flag <= 1'b1;
			end else begin
				out_result_97__flag<= 1'b0;
			end
			if(!(out_result_98__gfpga === out_result_98__bench) && !(out_result_98__bench === 1'bx)) begin
				out_result_98__flag <= 1'b1;
			end else begin
				out_result_98__flag<= 1'b0;
			end
			if(!(out_result_99__gfpga === out_result_99__bench) && !(out_result_99__bench === 1'bx)) begin
				out_result_99__flag <= 1'b1;
			end else begin
				out_result_99__flag<= 1'b0;
			end
			if(!(out_result_100__gfpga === out_result_100__bench) && !(out_result_100__bench === 1'bx)) begin
				out_result_100__flag <= 1'b1;
			end else begin
				out_result_100__flag<= 1'b0;
			end
			if(!(out_result_101__gfpga === out_result_101__bench) && !(out_result_101__bench === 1'bx)) begin
				out_result_101__flag <= 1'b1;
			end else begin
				out_result_101__flag<= 1'b0;
			end
			if(!(out_result_102__gfpga === out_result_102__bench) && !(out_result_102__bench === 1'bx)) begin
				out_result_102__flag <= 1'b1;
			end else begin
				out_result_102__flag<= 1'b0;
			end
			if(!(out_result_103__gfpga === out_result_103__bench) && !(out_result_103__bench === 1'bx)) begin
				out_result_103__flag <= 1'b1;
			end else begin
				out_result_103__flag<= 1'b0;
			end
			if(!(out_result_104__gfpga === out_result_104__bench) && !(out_result_104__bench === 1'bx)) begin
				out_result_104__flag <= 1'b1;
			end else begin
				out_result_104__flag<= 1'b0;
			end
			if(!(out_result_105__gfpga === out_result_105__bench) && !(out_result_105__bench === 1'bx)) begin
				out_result_105__flag <= 1'b1;
			end else begin
				out_result_105__flag<= 1'b0;
			end
			if(!(out_result_106__gfpga === out_result_106__bench) && !(out_result_106__bench === 1'bx)) begin
				out_result_106__flag <= 1'b1;
			end else begin
				out_result_106__flag<= 1'b0;
			end
			if(!(out_result_107__gfpga === out_result_107__bench) && !(out_result_107__bench === 1'bx)) begin
				out_result_107__flag <= 1'b1;
			end else begin
				out_result_107__flag<= 1'b0;
			end
			if(!(out_result_108__gfpga === out_result_108__bench) && !(out_result_108__bench === 1'bx)) begin
				out_result_108__flag <= 1'b1;
			end else begin
				out_result_108__flag<= 1'b0;
			end
			if(!(out_result_109__gfpga === out_result_109__bench) && !(out_result_109__bench === 1'bx)) begin
				out_result_109__flag <= 1'b1;
			end else begin
				out_result_109__flag<= 1'b0;
			end
			if(!(out_result_110__gfpga === out_result_110__bench) && !(out_result_110__bench === 1'bx)) begin
				out_result_110__flag <= 1'b1;
			end else begin
				out_result_110__flag<= 1'b0;
			end
			if(!(out_result_111__gfpga === out_result_111__bench) && !(out_result_111__bench === 1'bx)) begin
				out_result_111__flag <= 1'b1;
			end else begin
				out_result_111__flag<= 1'b0;
			end
			if(!(out_result_112__gfpga === out_result_112__bench) && !(out_result_112__bench === 1'bx)) begin
				out_result_112__flag <= 1'b1;
			end else begin
				out_result_112__flag<= 1'b0;
			end
			if(!(out_result_113__gfpga === out_result_113__bench) && !(out_result_113__bench === 1'bx)) begin
				out_result_113__flag <= 1'b1;
			end else begin
				out_result_113__flag<= 1'b0;
			end
			if(!(out_result_114__gfpga === out_result_114__bench) && !(out_result_114__bench === 1'bx)) begin
				out_result_114__flag <= 1'b1;
			end else begin
				out_result_114__flag<= 1'b0;
			end
			if(!(out_result_115__gfpga === out_result_115__bench) && !(out_result_115__bench === 1'bx)) begin
				out_result_115__flag <= 1'b1;
			end else begin
				out_result_115__flag<= 1'b0;
			end
			if(!(out_result_116__gfpga === out_result_116__bench) && !(out_result_116__bench === 1'bx)) begin
				out_result_116__flag <= 1'b1;
			end else begin
				out_result_116__flag<= 1'b0;
			end
			if(!(out_result_117__gfpga === out_result_117__bench) && !(out_result_117__bench === 1'bx)) begin
				out_result_117__flag <= 1'b1;
			end else begin
				out_result_117__flag<= 1'b0;
			end
			if(!(out_result_118__gfpga === out_result_118__bench) && !(out_result_118__bench === 1'bx)) begin
				out_result_118__flag <= 1'b1;
			end else begin
				out_result_118__flag<= 1'b0;
			end
			if(!(out_result_119__gfpga === out_result_119__bench) && !(out_result_119__bench === 1'bx)) begin
				out_result_119__flag <= 1'b1;
			end else begin
				out_result_119__flag<= 1'b0;
			end
			if(!(out_result_120__gfpga === out_result_120__bench) && !(out_result_120__bench === 1'bx)) begin
				out_result_120__flag <= 1'b1;
			end else begin
				out_result_120__flag<= 1'b0;
			end
			if(!(out_result_121__gfpga === out_result_121__bench) && !(out_result_121__bench === 1'bx)) begin
				out_result_121__flag <= 1'b1;
			end else begin
				out_result_121__flag<= 1'b0;
			end
			if(!(out_result_122__gfpga === out_result_122__bench) && !(out_result_122__bench === 1'bx)) begin
				out_result_122__flag <= 1'b1;
			end else begin
				out_result_122__flag<= 1'b0;
			end
			if(!(out_result_123__gfpga === out_result_123__bench) && !(out_result_123__bench === 1'bx)) begin
				out_result_123__flag <= 1'b1;
			end else begin
				out_result_123__flag<= 1'b0;
			end
			if(!(out_result_124__gfpga === out_result_124__bench) && !(out_result_124__bench === 1'bx)) begin
				out_result_124__flag <= 1'b1;
			end else begin
				out_result_124__flag<= 1'b0;
			end
			if(!(out_result_125__gfpga === out_result_125__bench) && !(out_result_125__bench === 1'bx)) begin
				out_result_125__flag <= 1'b1;
			end else begin
				out_result_125__flag<= 1'b0;
			end
			if(!(out_result_126__gfpga === out_result_126__bench) && !(out_result_126__bench === 1'bx)) begin
				out_result_126__flag <= 1'b1;
			end else begin
				out_result_126__flag<= 1'b0;
			end
			if(!(out_result_127__gfpga === out_result_127__bench) && !(out_result_127__bench === 1'bx)) begin
				out_result_127__flag <= 1'b1;
			end else begin
				out_result_127__flag<= 1'b0;
			end
		end
	end

	always@(posedge out_result_0__flag) begin
		if(out_result_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_1__flag) begin
		if(out_result_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_2__flag) begin
		if(out_result_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_3__flag) begin
		if(out_result_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_4__flag) begin
		if(out_result_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_5__flag) begin
		if(out_result_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_6__flag) begin
		if(out_result_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_7__flag) begin
		if(out_result_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_8__flag) begin
		if(out_result_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_9__flag) begin
		if(out_result_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_10__flag) begin
		if(out_result_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_11__flag) begin
		if(out_result_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_12__flag) begin
		if(out_result_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_13__flag) begin
		if(out_result_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_14__flag) begin
		if(out_result_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_15__flag) begin
		if(out_result_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_16__flag) begin
		if(out_result_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_17__flag) begin
		if(out_result_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_18__flag) begin
		if(out_result_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_19__flag) begin
		if(out_result_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_20__flag) begin
		if(out_result_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_21__flag) begin
		if(out_result_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_22__flag) begin
		if(out_result_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_23__flag) begin
		if(out_result_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_24__flag) begin
		if(out_result_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_25__flag) begin
		if(out_result_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_26__flag) begin
		if(out_result_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_27__flag) begin
		if(out_result_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_28__flag) begin
		if(out_result_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_29__flag) begin
		if(out_result_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_30__flag) begin
		if(out_result_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_31__flag) begin
		if(out_result_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_32__flag) begin
		if(out_result_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_33__flag) begin
		if(out_result_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_34__flag) begin
		if(out_result_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_35__flag) begin
		if(out_result_35__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_35__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_36__flag) begin
		if(out_result_36__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_36__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_37__flag) begin
		if(out_result_37__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_37__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_38__flag) begin
		if(out_result_38__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_38__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_39__flag) begin
		if(out_result_39__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_39__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_40__flag) begin
		if(out_result_40__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_40__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_41__flag) begin
		if(out_result_41__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_41__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_42__flag) begin
		if(out_result_42__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_42__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_43__flag) begin
		if(out_result_43__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_43__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_44__flag) begin
		if(out_result_44__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_44__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_45__flag) begin
		if(out_result_45__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_45__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_46__flag) begin
		if(out_result_46__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_46__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_47__flag) begin
		if(out_result_47__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_47__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_48__flag) begin
		if(out_result_48__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_48__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_49__flag) begin
		if(out_result_49__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_49__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_50__flag) begin
		if(out_result_50__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_50__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_51__flag) begin
		if(out_result_51__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_51__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_52__flag) begin
		if(out_result_52__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_52__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_53__flag) begin
		if(out_result_53__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_53__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_54__flag) begin
		if(out_result_54__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_54__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_55__flag) begin
		if(out_result_55__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_55__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_56__flag) begin
		if(out_result_56__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_56__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_57__flag) begin
		if(out_result_57__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_57__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_58__flag) begin
		if(out_result_58__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_58__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_59__flag) begin
		if(out_result_59__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_59__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_60__flag) begin
		if(out_result_60__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_60__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_61__flag) begin
		if(out_result_61__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_61__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_62__flag) begin
		if(out_result_62__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_62__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_63__flag) begin
		if(out_result_63__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_63__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_64__flag) begin
		if(out_result_64__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_64__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_65__flag) begin
		if(out_result_65__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_65__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_66__flag) begin
		if(out_result_66__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_66__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_67__flag) begin
		if(out_result_67__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_67__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_68__flag) begin
		if(out_result_68__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_68__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_69__flag) begin
		if(out_result_69__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_69__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_70__flag) begin
		if(out_result_70__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_70__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_71__flag) begin
		if(out_result_71__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_71__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_72__flag) begin
		if(out_result_72__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_72__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_73__flag) begin
		if(out_result_73__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_73__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_74__flag) begin
		if(out_result_74__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_74__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_75__flag) begin
		if(out_result_75__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_75__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_76__flag) begin
		if(out_result_76__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_76__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_77__flag) begin
		if(out_result_77__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_77__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_78__flag) begin
		if(out_result_78__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_78__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_79__flag) begin
		if(out_result_79__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_79__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_80__flag) begin
		if(out_result_80__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_80__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_81__flag) begin
		if(out_result_81__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_81__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_82__flag) begin
		if(out_result_82__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_82__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_83__flag) begin
		if(out_result_83__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_83__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_84__flag) begin
		if(out_result_84__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_84__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_85__flag) begin
		if(out_result_85__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_85__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_86__flag) begin
		if(out_result_86__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_86__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_87__flag) begin
		if(out_result_87__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_87__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_88__flag) begin
		if(out_result_88__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_88__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_89__flag) begin
		if(out_result_89__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_89__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_90__flag) begin
		if(out_result_90__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_90__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_91__flag) begin
		if(out_result_91__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_91__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_92__flag) begin
		if(out_result_92__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_92__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_93__flag) begin
		if(out_result_93__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_93__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_94__flag) begin
		if(out_result_94__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_94__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_95__flag) begin
		if(out_result_95__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_95__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_96__flag) begin
		if(out_result_96__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_96__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_97__flag) begin
		if(out_result_97__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_97__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_98__flag) begin
		if(out_result_98__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_98__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_99__flag) begin
		if(out_result_99__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_99__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_100__flag) begin
		if(out_result_100__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_100__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_101__flag) begin
		if(out_result_101__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_101__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_102__flag) begin
		if(out_result_102__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_102__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_103__flag) begin
		if(out_result_103__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_103__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_104__flag) begin
		if(out_result_104__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_104__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_105__flag) begin
		if(out_result_105__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_105__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_106__flag) begin
		if(out_result_106__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_106__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_107__flag) begin
		if(out_result_107__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_107__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_108__flag) begin
		if(out_result_108__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_108__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_109__flag) begin
		if(out_result_109__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_109__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_110__flag) begin
		if(out_result_110__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_110__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_111__flag) begin
		if(out_result_111__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_111__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_112__flag) begin
		if(out_result_112__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_112__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_113__flag) begin
		if(out_result_113__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_113__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_114__flag) begin
		if(out_result_114__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_114__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_115__flag) begin
		if(out_result_115__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_115__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_116__flag) begin
		if(out_result_116__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_116__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_117__flag) begin
		if(out_result_117__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_117__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_118__flag) begin
		if(out_result_118__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_118__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_119__flag) begin
		if(out_result_119__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_119__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_120__flag) begin
		if(out_result_120__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_120__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_121__flag) begin
		if(out_result_121__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_121__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_122__flag) begin
		if(out_result_122__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_122__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_123__flag) begin
		if(out_result_123__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_123__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_124__flag) begin
		if(out_result_124__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_124__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_125__flag) begin
		if(out_result_125__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_125__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_126__flag) begin
		if(out_result_126__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_126__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge out_result_127__flag) begin
		if(out_result_127__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_result_127__gfpga at time = %t", $realtime);
		end
	end


// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("counter_formal.vcd");
		$dumpvars(1, counter_top_formal_verification_random_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#20
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for counter_top_formal_verification_random_tb -----

//----- Default net type -----
// `default_nettype none

