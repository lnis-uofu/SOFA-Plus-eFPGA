

module fpga_top
(
  input [0:0] config_enable,
  input [0:0] pReset,
  input [0:0] prog_clk,
  input [0:0] Test_en,
  input [0:0] IO_ISOL_N,
  input [0:0] clk,
  input [0:0] reset,
  input [0:143] gfpga_pad_sofa_plus_io_SOC_IN,
  output [0:143] gfpga_pad_sofa_plus_io_SOC_OUT,
  output [0:143] gfpga_pad_sofa_plus_io_SOC_DIR,
  input [0:11] ccff_head,
  output [0:11] ccff_tail
);

  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_ccff_tail;
  wire [0:19] cbx_1__0__0_chanx_left_out;
  wire [0:19] cbx_1__0__0_chanx_right_out;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_ccff_tail;
  wire [0:19] cbx_1__0__10_chanx_left_out;
  wire [0:19] cbx_1__0__10_chanx_right_out;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_ccff_tail;
  wire [0:19] cbx_1__0__11_chanx_left_out;
  wire [0:19] cbx_1__0__11_chanx_right_out;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_ccff_tail;
  wire [0:19] cbx_1__0__1_chanx_left_out;
  wire [0:19] cbx_1__0__1_chanx_right_out;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_ccff_tail;
  wire [0:19] cbx_1__0__2_chanx_left_out;
  wire [0:19] cbx_1__0__2_chanx_right_out;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_ccff_tail;
  wire [0:19] cbx_1__0__3_chanx_left_out;
  wire [0:19] cbx_1__0__3_chanx_right_out;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_ccff_tail;
  wire [0:19] cbx_1__0__4_chanx_left_out;
  wire [0:19] cbx_1__0__4_chanx_right_out;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_ccff_tail;
  wire [0:19] cbx_1__0__5_chanx_left_out;
  wire [0:19] cbx_1__0__5_chanx_right_out;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_ccff_tail;
  wire [0:19] cbx_1__0__6_chanx_left_out;
  wire [0:19] cbx_1__0__6_chanx_right_out;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_ccff_tail;
  wire [0:19] cbx_1__0__7_chanx_left_out;
  wire [0:19] cbx_1__0__7_chanx_right_out;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_ccff_tail;
  wire [0:19] cbx_1__0__8_chanx_left_out;
  wire [0:19] cbx_1__0__8_chanx_right_out;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_ccff_tail;
  wire [0:19] cbx_1__0__9_chanx_left_out;
  wire [0:19] cbx_1__0__9_chanx_right_out;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__0_ccff_tail;
  wire [0:19] cbx_1__12__0_chanx_left_out;
  wire [0:19] cbx_1__12__0_chanx_right_out;
  wire [0:0] cbx_1__12__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__10_ccff_tail;
  wire [0:19] cbx_1__12__10_chanx_left_out;
  wire [0:19] cbx_1__12__10_chanx_right_out;
  wire [0:0] cbx_1__12__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__11_ccff_tail;
  wire [0:19] cbx_1__12__11_chanx_left_out;
  wire [0:19] cbx_1__12__11_chanx_right_out;
  wire [0:0] cbx_1__12__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__1_ccff_tail;
  wire [0:19] cbx_1__12__1_chanx_left_out;
  wire [0:19] cbx_1__12__1_chanx_right_out;
  wire [0:0] cbx_1__12__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__2_ccff_tail;
  wire [0:19] cbx_1__12__2_chanx_left_out;
  wire [0:19] cbx_1__12__2_chanx_right_out;
  wire [0:0] cbx_1__12__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__3_ccff_tail;
  wire [0:19] cbx_1__12__3_chanx_left_out;
  wire [0:19] cbx_1__12__3_chanx_right_out;
  wire [0:0] cbx_1__12__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__4_ccff_tail;
  wire [0:19] cbx_1__12__4_chanx_left_out;
  wire [0:19] cbx_1__12__4_chanx_right_out;
  wire [0:0] cbx_1__12__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__5_ccff_tail;
  wire [0:19] cbx_1__12__5_chanx_left_out;
  wire [0:19] cbx_1__12__5_chanx_right_out;
  wire [0:0] cbx_1__12__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__6_ccff_tail;
  wire [0:19] cbx_1__12__6_chanx_left_out;
  wire [0:19] cbx_1__12__6_chanx_right_out;
  wire [0:0] cbx_1__12__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__7_ccff_tail;
  wire [0:19] cbx_1__12__7_chanx_left_out;
  wire [0:19] cbx_1__12__7_chanx_right_out;
  wire [0:0] cbx_1__12__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__8_ccff_tail;
  wire [0:19] cbx_1__12__8_chanx_left_out;
  wire [0:19] cbx_1__12__8_chanx_right_out;
  wire [0:0] cbx_1__12__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__9_ccff_tail;
  wire [0:19] cbx_1__12__9_chanx_left_out;
  wire [0:19] cbx_1__12__9_chanx_right_out;
  wire [0:0] cbx_1__12__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__0_ccff_tail;
  wire [0:19] cbx_1__1__0_chanx_left_out;
  wire [0:19] cbx_1__1__0_chanx_right_out;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__100_ccff_tail;
  wire [0:19] cbx_1__1__100_chanx_left_out;
  wire [0:19] cbx_1__1__100_chanx_right_out;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__101_ccff_tail;
  wire [0:19] cbx_1__1__101_chanx_left_out;
  wire [0:19] cbx_1__1__101_chanx_right_out;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__102_ccff_tail;
  wire [0:19] cbx_1__1__102_chanx_left_out;
  wire [0:19] cbx_1__1__102_chanx_right_out;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__103_ccff_tail;
  wire [0:19] cbx_1__1__103_chanx_left_out;
  wire [0:19] cbx_1__1__103_chanx_right_out;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__104_ccff_tail;
  wire [0:19] cbx_1__1__104_chanx_left_out;
  wire [0:19] cbx_1__1__104_chanx_right_out;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__105_ccff_tail;
  wire [0:19] cbx_1__1__105_chanx_left_out;
  wire [0:19] cbx_1__1__105_chanx_right_out;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__106_ccff_tail;
  wire [0:19] cbx_1__1__106_chanx_left_out;
  wire [0:19] cbx_1__1__106_chanx_right_out;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__107_ccff_tail;
  wire [0:19] cbx_1__1__107_chanx_left_out;
  wire [0:19] cbx_1__1__107_chanx_right_out;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__10_ccff_tail;
  wire [0:19] cbx_1__1__10_chanx_left_out;
  wire [0:19] cbx_1__1__10_chanx_right_out;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__11_ccff_tail;
  wire [0:19] cbx_1__1__11_chanx_left_out;
  wire [0:19] cbx_1__1__11_chanx_right_out;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__12_ccff_tail;
  wire [0:19] cbx_1__1__12_chanx_left_out;
  wire [0:19] cbx_1__1__12_chanx_right_out;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__13_ccff_tail;
  wire [0:19] cbx_1__1__13_chanx_left_out;
  wire [0:19] cbx_1__1__13_chanx_right_out;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__14_ccff_tail;
  wire [0:19] cbx_1__1__14_chanx_left_out;
  wire [0:19] cbx_1__1__14_chanx_right_out;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__15_ccff_tail;
  wire [0:19] cbx_1__1__15_chanx_left_out;
  wire [0:19] cbx_1__1__15_chanx_right_out;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__16_ccff_tail;
  wire [0:19] cbx_1__1__16_chanx_left_out;
  wire [0:19] cbx_1__1__16_chanx_right_out;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__17_ccff_tail;
  wire [0:19] cbx_1__1__17_chanx_left_out;
  wire [0:19] cbx_1__1__17_chanx_right_out;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__18_ccff_tail;
  wire [0:19] cbx_1__1__18_chanx_left_out;
  wire [0:19] cbx_1__1__18_chanx_right_out;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__19_ccff_tail;
  wire [0:19] cbx_1__1__19_chanx_left_out;
  wire [0:19] cbx_1__1__19_chanx_right_out;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__1_ccff_tail;
  wire [0:19] cbx_1__1__1_chanx_left_out;
  wire [0:19] cbx_1__1__1_chanx_right_out;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__20_ccff_tail;
  wire [0:19] cbx_1__1__20_chanx_left_out;
  wire [0:19] cbx_1__1__20_chanx_right_out;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__21_ccff_tail;
  wire [0:19] cbx_1__1__21_chanx_left_out;
  wire [0:19] cbx_1__1__21_chanx_right_out;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__22_ccff_tail;
  wire [0:19] cbx_1__1__22_chanx_left_out;
  wire [0:19] cbx_1__1__22_chanx_right_out;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__23_ccff_tail;
  wire [0:19] cbx_1__1__23_chanx_left_out;
  wire [0:19] cbx_1__1__23_chanx_right_out;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__24_ccff_tail;
  wire [0:19] cbx_1__1__24_chanx_left_out;
  wire [0:19] cbx_1__1__24_chanx_right_out;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__25_ccff_tail;
  wire [0:19] cbx_1__1__25_chanx_left_out;
  wire [0:19] cbx_1__1__25_chanx_right_out;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__26_ccff_tail;
  wire [0:19] cbx_1__1__26_chanx_left_out;
  wire [0:19] cbx_1__1__26_chanx_right_out;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__27_ccff_tail;
  wire [0:19] cbx_1__1__27_chanx_left_out;
  wire [0:19] cbx_1__1__27_chanx_right_out;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__28_ccff_tail;
  wire [0:19] cbx_1__1__28_chanx_left_out;
  wire [0:19] cbx_1__1__28_chanx_right_out;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__29_ccff_tail;
  wire [0:19] cbx_1__1__29_chanx_left_out;
  wire [0:19] cbx_1__1__29_chanx_right_out;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__2_ccff_tail;
  wire [0:19] cbx_1__1__2_chanx_left_out;
  wire [0:19] cbx_1__1__2_chanx_right_out;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__30_ccff_tail;
  wire [0:19] cbx_1__1__30_chanx_left_out;
  wire [0:19] cbx_1__1__30_chanx_right_out;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__31_ccff_tail;
  wire [0:19] cbx_1__1__31_chanx_left_out;
  wire [0:19] cbx_1__1__31_chanx_right_out;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__32_ccff_tail;
  wire [0:19] cbx_1__1__32_chanx_left_out;
  wire [0:19] cbx_1__1__32_chanx_right_out;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__33_ccff_tail;
  wire [0:19] cbx_1__1__33_chanx_left_out;
  wire [0:19] cbx_1__1__33_chanx_right_out;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__34_ccff_tail;
  wire [0:19] cbx_1__1__34_chanx_left_out;
  wire [0:19] cbx_1__1__34_chanx_right_out;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__35_ccff_tail;
  wire [0:19] cbx_1__1__35_chanx_left_out;
  wire [0:19] cbx_1__1__35_chanx_right_out;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__36_ccff_tail;
  wire [0:19] cbx_1__1__36_chanx_left_out;
  wire [0:19] cbx_1__1__36_chanx_right_out;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__37_ccff_tail;
  wire [0:19] cbx_1__1__37_chanx_left_out;
  wire [0:19] cbx_1__1__37_chanx_right_out;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__38_ccff_tail;
  wire [0:19] cbx_1__1__38_chanx_left_out;
  wire [0:19] cbx_1__1__38_chanx_right_out;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__39_ccff_tail;
  wire [0:19] cbx_1__1__39_chanx_left_out;
  wire [0:19] cbx_1__1__39_chanx_right_out;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__3_ccff_tail;
  wire [0:19] cbx_1__1__3_chanx_left_out;
  wire [0:19] cbx_1__1__3_chanx_right_out;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__40_ccff_tail;
  wire [0:19] cbx_1__1__40_chanx_left_out;
  wire [0:19] cbx_1__1__40_chanx_right_out;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__41_ccff_tail;
  wire [0:19] cbx_1__1__41_chanx_left_out;
  wire [0:19] cbx_1__1__41_chanx_right_out;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__42_ccff_tail;
  wire [0:19] cbx_1__1__42_chanx_left_out;
  wire [0:19] cbx_1__1__42_chanx_right_out;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__43_ccff_tail;
  wire [0:19] cbx_1__1__43_chanx_left_out;
  wire [0:19] cbx_1__1__43_chanx_right_out;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__44_ccff_tail;
  wire [0:19] cbx_1__1__44_chanx_left_out;
  wire [0:19] cbx_1__1__44_chanx_right_out;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__45_ccff_tail;
  wire [0:19] cbx_1__1__45_chanx_left_out;
  wire [0:19] cbx_1__1__45_chanx_right_out;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__46_ccff_tail;
  wire [0:19] cbx_1__1__46_chanx_left_out;
  wire [0:19] cbx_1__1__46_chanx_right_out;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__47_ccff_tail;
  wire [0:19] cbx_1__1__47_chanx_left_out;
  wire [0:19] cbx_1__1__47_chanx_right_out;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__48_ccff_tail;
  wire [0:19] cbx_1__1__48_chanx_left_out;
  wire [0:19] cbx_1__1__48_chanx_right_out;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__49_ccff_tail;
  wire [0:19] cbx_1__1__49_chanx_left_out;
  wire [0:19] cbx_1__1__49_chanx_right_out;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__4_ccff_tail;
  wire [0:19] cbx_1__1__4_chanx_left_out;
  wire [0:19] cbx_1__1__4_chanx_right_out;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__50_ccff_tail;
  wire [0:19] cbx_1__1__50_chanx_left_out;
  wire [0:19] cbx_1__1__50_chanx_right_out;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__51_ccff_tail;
  wire [0:19] cbx_1__1__51_chanx_left_out;
  wire [0:19] cbx_1__1__51_chanx_right_out;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__52_ccff_tail;
  wire [0:19] cbx_1__1__52_chanx_left_out;
  wire [0:19] cbx_1__1__52_chanx_right_out;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__53_ccff_tail;
  wire [0:19] cbx_1__1__53_chanx_left_out;
  wire [0:19] cbx_1__1__53_chanx_right_out;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__54_ccff_tail;
  wire [0:19] cbx_1__1__54_chanx_left_out;
  wire [0:19] cbx_1__1__54_chanx_right_out;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__55_ccff_tail;
  wire [0:19] cbx_1__1__55_chanx_left_out;
  wire [0:19] cbx_1__1__55_chanx_right_out;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__56_ccff_tail;
  wire [0:19] cbx_1__1__56_chanx_left_out;
  wire [0:19] cbx_1__1__56_chanx_right_out;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__57_ccff_tail;
  wire [0:19] cbx_1__1__57_chanx_left_out;
  wire [0:19] cbx_1__1__57_chanx_right_out;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__58_ccff_tail;
  wire [0:19] cbx_1__1__58_chanx_left_out;
  wire [0:19] cbx_1__1__58_chanx_right_out;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__59_ccff_tail;
  wire [0:19] cbx_1__1__59_chanx_left_out;
  wire [0:19] cbx_1__1__59_chanx_right_out;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__5_ccff_tail;
  wire [0:19] cbx_1__1__5_chanx_left_out;
  wire [0:19] cbx_1__1__5_chanx_right_out;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__60_ccff_tail;
  wire [0:19] cbx_1__1__60_chanx_left_out;
  wire [0:19] cbx_1__1__60_chanx_right_out;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__61_ccff_tail;
  wire [0:19] cbx_1__1__61_chanx_left_out;
  wire [0:19] cbx_1__1__61_chanx_right_out;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__62_ccff_tail;
  wire [0:19] cbx_1__1__62_chanx_left_out;
  wire [0:19] cbx_1__1__62_chanx_right_out;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__63_ccff_tail;
  wire [0:19] cbx_1__1__63_chanx_left_out;
  wire [0:19] cbx_1__1__63_chanx_right_out;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__64_ccff_tail;
  wire [0:19] cbx_1__1__64_chanx_left_out;
  wire [0:19] cbx_1__1__64_chanx_right_out;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__65_ccff_tail;
  wire [0:19] cbx_1__1__65_chanx_left_out;
  wire [0:19] cbx_1__1__65_chanx_right_out;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__66_ccff_tail;
  wire [0:19] cbx_1__1__66_chanx_left_out;
  wire [0:19] cbx_1__1__66_chanx_right_out;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__67_ccff_tail;
  wire [0:19] cbx_1__1__67_chanx_left_out;
  wire [0:19] cbx_1__1__67_chanx_right_out;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__68_ccff_tail;
  wire [0:19] cbx_1__1__68_chanx_left_out;
  wire [0:19] cbx_1__1__68_chanx_right_out;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__69_ccff_tail;
  wire [0:19] cbx_1__1__69_chanx_left_out;
  wire [0:19] cbx_1__1__69_chanx_right_out;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__6_ccff_tail;
  wire [0:19] cbx_1__1__6_chanx_left_out;
  wire [0:19] cbx_1__1__6_chanx_right_out;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__70_ccff_tail;
  wire [0:19] cbx_1__1__70_chanx_left_out;
  wire [0:19] cbx_1__1__70_chanx_right_out;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__71_ccff_tail;
  wire [0:19] cbx_1__1__71_chanx_left_out;
  wire [0:19] cbx_1__1__71_chanx_right_out;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__72_ccff_tail;
  wire [0:19] cbx_1__1__72_chanx_left_out;
  wire [0:19] cbx_1__1__72_chanx_right_out;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__73_ccff_tail;
  wire [0:19] cbx_1__1__73_chanx_left_out;
  wire [0:19] cbx_1__1__73_chanx_right_out;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__74_ccff_tail;
  wire [0:19] cbx_1__1__74_chanx_left_out;
  wire [0:19] cbx_1__1__74_chanx_right_out;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__75_ccff_tail;
  wire [0:19] cbx_1__1__75_chanx_left_out;
  wire [0:19] cbx_1__1__75_chanx_right_out;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__76_ccff_tail;
  wire [0:19] cbx_1__1__76_chanx_left_out;
  wire [0:19] cbx_1__1__76_chanx_right_out;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__77_ccff_tail;
  wire [0:19] cbx_1__1__77_chanx_left_out;
  wire [0:19] cbx_1__1__77_chanx_right_out;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__78_ccff_tail;
  wire [0:19] cbx_1__1__78_chanx_left_out;
  wire [0:19] cbx_1__1__78_chanx_right_out;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__79_ccff_tail;
  wire [0:19] cbx_1__1__79_chanx_left_out;
  wire [0:19] cbx_1__1__79_chanx_right_out;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__7_ccff_tail;
  wire [0:19] cbx_1__1__7_chanx_left_out;
  wire [0:19] cbx_1__1__7_chanx_right_out;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__80_ccff_tail;
  wire [0:19] cbx_1__1__80_chanx_left_out;
  wire [0:19] cbx_1__1__80_chanx_right_out;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__81_ccff_tail;
  wire [0:19] cbx_1__1__81_chanx_left_out;
  wire [0:19] cbx_1__1__81_chanx_right_out;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__82_ccff_tail;
  wire [0:19] cbx_1__1__82_chanx_left_out;
  wire [0:19] cbx_1__1__82_chanx_right_out;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__83_ccff_tail;
  wire [0:19] cbx_1__1__83_chanx_left_out;
  wire [0:19] cbx_1__1__83_chanx_right_out;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__84_ccff_tail;
  wire [0:19] cbx_1__1__84_chanx_left_out;
  wire [0:19] cbx_1__1__84_chanx_right_out;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__85_ccff_tail;
  wire [0:19] cbx_1__1__85_chanx_left_out;
  wire [0:19] cbx_1__1__85_chanx_right_out;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__86_ccff_tail;
  wire [0:19] cbx_1__1__86_chanx_left_out;
  wire [0:19] cbx_1__1__86_chanx_right_out;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__87_ccff_tail;
  wire [0:19] cbx_1__1__87_chanx_left_out;
  wire [0:19] cbx_1__1__87_chanx_right_out;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__88_ccff_tail;
  wire [0:19] cbx_1__1__88_chanx_left_out;
  wire [0:19] cbx_1__1__88_chanx_right_out;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__89_ccff_tail;
  wire [0:19] cbx_1__1__89_chanx_left_out;
  wire [0:19] cbx_1__1__89_chanx_right_out;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__8_ccff_tail;
  wire [0:19] cbx_1__1__8_chanx_left_out;
  wire [0:19] cbx_1__1__8_chanx_right_out;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__90_ccff_tail;
  wire [0:19] cbx_1__1__90_chanx_left_out;
  wire [0:19] cbx_1__1__90_chanx_right_out;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__91_ccff_tail;
  wire [0:19] cbx_1__1__91_chanx_left_out;
  wire [0:19] cbx_1__1__91_chanx_right_out;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__92_ccff_tail;
  wire [0:19] cbx_1__1__92_chanx_left_out;
  wire [0:19] cbx_1__1__92_chanx_right_out;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__93_ccff_tail;
  wire [0:19] cbx_1__1__93_chanx_left_out;
  wire [0:19] cbx_1__1__93_chanx_right_out;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__94_ccff_tail;
  wire [0:19] cbx_1__1__94_chanx_left_out;
  wire [0:19] cbx_1__1__94_chanx_right_out;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__95_ccff_tail;
  wire [0:19] cbx_1__1__95_chanx_left_out;
  wire [0:19] cbx_1__1__95_chanx_right_out;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__96_ccff_tail;
  wire [0:19] cbx_1__1__96_chanx_left_out;
  wire [0:19] cbx_1__1__96_chanx_right_out;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__97_ccff_tail;
  wire [0:19] cbx_1__1__97_chanx_left_out;
  wire [0:19] cbx_1__1__97_chanx_right_out;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__98_ccff_tail;
  wire [0:19] cbx_1__1__98_chanx_left_out;
  wire [0:19] cbx_1__1__98_chanx_right_out;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__99_ccff_tail;
  wire [0:19] cbx_1__1__99_chanx_left_out;
  wire [0:19] cbx_1__1__99_chanx_right_out;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__9_ccff_tail;
  wire [0:19] cbx_1__1__9_chanx_left_out;
  wire [0:19] cbx_1__1__9_chanx_right_out;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__0_ccff_tail;
  wire [0:19] cbx_1__3__0_chanx_left_out;
  wire [0:19] cbx_1__3__0_chanx_right_out;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__10_ccff_tail;
  wire [0:19] cbx_1__3__10_chanx_left_out;
  wire [0:19] cbx_1__3__10_chanx_right_out;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__11_ccff_tail;
  wire [0:19] cbx_1__3__11_chanx_left_out;
  wire [0:19] cbx_1__3__11_chanx_right_out;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__1_ccff_tail;
  wire [0:19] cbx_1__3__1_chanx_left_out;
  wire [0:19] cbx_1__3__1_chanx_right_out;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__2_ccff_tail;
  wire [0:19] cbx_1__3__2_chanx_left_out;
  wire [0:19] cbx_1__3__2_chanx_right_out;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__3_ccff_tail;
  wire [0:19] cbx_1__3__3_chanx_left_out;
  wire [0:19] cbx_1__3__3_chanx_right_out;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__4_ccff_tail;
  wire [0:19] cbx_1__3__4_chanx_left_out;
  wire [0:19] cbx_1__3__4_chanx_right_out;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__5_ccff_tail;
  wire [0:19] cbx_1__3__5_chanx_left_out;
  wire [0:19] cbx_1__3__5_chanx_right_out;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__6_ccff_tail;
  wire [0:19] cbx_1__3__6_chanx_left_out;
  wire [0:19] cbx_1__3__6_chanx_right_out;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__7_ccff_tail;
  wire [0:19] cbx_1__3__7_chanx_left_out;
  wire [0:19] cbx_1__3__7_chanx_right_out;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__8_ccff_tail;
  wire [0:19] cbx_1__3__8_chanx_left_out;
  wire [0:19] cbx_1__3__8_chanx_right_out;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__9_ccff_tail;
  wire [0:19] cbx_1__3__9_chanx_left_out;
  wire [0:19] cbx_1__3__9_chanx_right_out;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__0_ccff_tail;
  wire [0:19] cbx_2__3__0_chanx_left_out;
  wire [0:19] cbx_2__3__0_chanx_right_out;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__10_ccff_tail;
  wire [0:19] cbx_2__3__10_chanx_left_out;
  wire [0:19] cbx_2__3__10_chanx_right_out;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__11_ccff_tail;
  wire [0:19] cbx_2__3__11_chanx_left_out;
  wire [0:19] cbx_2__3__11_chanx_right_out;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__1_ccff_tail;
  wire [0:19] cbx_2__3__1_chanx_left_out;
  wire [0:19] cbx_2__3__1_chanx_right_out;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__2_ccff_tail;
  wire [0:19] cbx_2__3__2_chanx_left_out;
  wire [0:19] cbx_2__3__2_chanx_right_out;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__3_ccff_tail;
  wire [0:19] cbx_2__3__3_chanx_left_out;
  wire [0:19] cbx_2__3__3_chanx_right_out;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__4_ccff_tail;
  wire [0:19] cbx_2__3__4_chanx_left_out;
  wire [0:19] cbx_2__3__4_chanx_right_out;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__5_ccff_tail;
  wire [0:19] cbx_2__3__5_chanx_left_out;
  wire [0:19] cbx_2__3__5_chanx_right_out;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__6_ccff_tail;
  wire [0:19] cbx_2__3__6_chanx_left_out;
  wire [0:19] cbx_2__3__6_chanx_right_out;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__7_ccff_tail;
  wire [0:19] cbx_2__3__7_chanx_left_out;
  wire [0:19] cbx_2__3__7_chanx_right_out;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__8_ccff_tail;
  wire [0:19] cbx_2__3__8_chanx_left_out;
  wire [0:19] cbx_2__3__8_chanx_right_out;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__9_ccff_tail;
  wire [0:19] cbx_2__3__9_chanx_left_out;
  wire [0:19] cbx_2__3__9_chanx_right_out;
  wire [0:0] cby_0__1__0_ccff_tail;
  wire [0:19] cby_0__1__0_chany_bottom_out;
  wire [0:19] cby_0__1__0_chany_top_out;
  wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__10_ccff_tail;
  wire [0:19] cby_0__1__10_chany_bottom_out;
  wire [0:19] cby_0__1__10_chany_top_out;
  wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__11_ccff_tail;
  wire [0:19] cby_0__1__11_chany_bottom_out;
  wire [0:19] cby_0__1__11_chany_top_out;
  wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__1_ccff_tail;
  wire [0:19] cby_0__1__1_chany_bottom_out;
  wire [0:19] cby_0__1__1_chany_top_out;
  wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__2_ccff_tail;
  wire [0:19] cby_0__1__2_chany_bottom_out;
  wire [0:19] cby_0__1__2_chany_top_out;
  wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__3_ccff_tail;
  wire [0:19] cby_0__1__3_chany_bottom_out;
  wire [0:19] cby_0__1__3_chany_top_out;
  wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__4_ccff_tail;
  wire [0:19] cby_0__1__4_chany_bottom_out;
  wire [0:19] cby_0__1__4_chany_top_out;
  wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__5_ccff_tail;
  wire [0:19] cby_0__1__5_chany_bottom_out;
  wire [0:19] cby_0__1__5_chany_top_out;
  wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__6_ccff_tail;
  wire [0:19] cby_0__1__6_chany_bottom_out;
  wire [0:19] cby_0__1__6_chany_top_out;
  wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__7_ccff_tail;
  wire [0:19] cby_0__1__7_chany_bottom_out;
  wire [0:19] cby_0__1__7_chany_top_out;
  wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__8_ccff_tail;
  wire [0:19] cby_0__1__8_chany_bottom_out;
  wire [0:19] cby_0__1__8_chany_top_out;
  wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__9_ccff_tail;
  wire [0:19] cby_0__1__9_chany_bottom_out;
  wire [0:19] cby_0__1__9_chany_top_out;
  wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__0_ccff_tail;
  wire [0:19] cby_12__1__0_chany_bottom_out;
  wire [0:19] cby_12__1__0_chany_top_out;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__1_ccff_tail;
  wire [0:19] cby_12__1__1_chany_bottom_out;
  wire [0:19] cby_12__1__1_chany_top_out;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__2_ccff_tail;
  wire [0:19] cby_12__1__2_chany_bottom_out;
  wire [0:19] cby_12__1__2_chany_top_out;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__3_ccff_tail;
  wire [0:19] cby_12__1__3_chany_bottom_out;
  wire [0:19] cby_12__1__3_chany_top_out;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__4_ccff_tail;
  wire [0:19] cby_12__1__4_chany_bottom_out;
  wire [0:19] cby_12__1__4_chany_top_out;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__5_ccff_tail;
  wire [0:19] cby_12__1__5_chany_bottom_out;
  wire [0:19] cby_12__1__5_chany_top_out;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__6_ccff_tail;
  wire [0:19] cby_12__1__6_chany_bottom_out;
  wire [0:19] cby_12__1__6_chany_top_out;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__7_ccff_tail;
  wire [0:19] cby_12__1__7_chany_bottom_out;
  wire [0:19] cby_12__1__7_chany_top_out;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__8_ccff_tail;
  wire [0:19] cby_12__1__8_chany_bottom_out;
  wire [0:19] cby_12__1__8_chany_top_out;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__9_ccff_tail;
  wire [0:19] cby_12__1__9_chany_bottom_out;
  wire [0:19] cby_12__1__9_chany_top_out;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__3__0_ccff_tail;
  wire [0:19] cby_12__3__0_chany_bottom_out;
  wire [0:19] cby_12__3__0_chany_top_out;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_12__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__3__1_ccff_tail;
  wire [0:19] cby_12__3__1_chany_bottom_out;
  wire [0:19] cby_12__3__1_chany_top_out;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_12__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_1__1__0_ccff_tail;
  wire [0:19] cby_1__1__0_chany_bottom_out;
  wire [0:19] cby_1__1__0_chany_top_out;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__100_ccff_tail;
  wire [0:19] cby_1__1__100_chany_bottom_out;
  wire [0:19] cby_1__1__100_chany_top_out;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__101_ccff_tail;
  wire [0:19] cby_1__1__101_chany_bottom_out;
  wire [0:19] cby_1__1__101_chany_top_out;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__102_ccff_tail;
  wire [0:19] cby_1__1__102_chany_bottom_out;
  wire [0:19] cby_1__1__102_chany_top_out;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__103_ccff_tail;
  wire [0:19] cby_1__1__103_chany_bottom_out;
  wire [0:19] cby_1__1__103_chany_top_out;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__104_ccff_tail;
  wire [0:19] cby_1__1__104_chany_bottom_out;
  wire [0:19] cby_1__1__104_chany_top_out;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__105_ccff_tail;
  wire [0:19] cby_1__1__105_chany_bottom_out;
  wire [0:19] cby_1__1__105_chany_top_out;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__106_ccff_tail;
  wire [0:19] cby_1__1__106_chany_bottom_out;
  wire [0:19] cby_1__1__106_chany_top_out;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__107_ccff_tail;
  wire [0:19] cby_1__1__107_chany_bottom_out;
  wire [0:19] cby_1__1__107_chany_top_out;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__108_ccff_tail;
  wire [0:19] cby_1__1__108_chany_bottom_out;
  wire [0:19] cby_1__1__108_chany_top_out;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__109_ccff_tail;
  wire [0:19] cby_1__1__109_chany_bottom_out;
  wire [0:19] cby_1__1__109_chany_top_out;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__10_ccff_tail;
  wire [0:19] cby_1__1__10_chany_bottom_out;
  wire [0:19] cby_1__1__10_chany_top_out;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__11_ccff_tail;
  wire [0:19] cby_1__1__11_chany_bottom_out;
  wire [0:19] cby_1__1__11_chany_top_out;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__12_ccff_tail;
  wire [0:19] cby_1__1__12_chany_bottom_out;
  wire [0:19] cby_1__1__12_chany_top_out;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__13_ccff_tail;
  wire [0:19] cby_1__1__13_chany_bottom_out;
  wire [0:19] cby_1__1__13_chany_top_out;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__14_ccff_tail;
  wire [0:19] cby_1__1__14_chany_bottom_out;
  wire [0:19] cby_1__1__14_chany_top_out;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__15_ccff_tail;
  wire [0:19] cby_1__1__15_chany_bottom_out;
  wire [0:19] cby_1__1__15_chany_top_out;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__16_ccff_tail;
  wire [0:19] cby_1__1__16_chany_bottom_out;
  wire [0:19] cby_1__1__16_chany_top_out;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__17_ccff_tail;
  wire [0:19] cby_1__1__17_chany_bottom_out;
  wire [0:19] cby_1__1__17_chany_top_out;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__18_ccff_tail;
  wire [0:19] cby_1__1__18_chany_bottom_out;
  wire [0:19] cby_1__1__18_chany_top_out;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__19_ccff_tail;
  wire [0:19] cby_1__1__19_chany_bottom_out;
  wire [0:19] cby_1__1__19_chany_top_out;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__1_ccff_tail;
  wire [0:19] cby_1__1__1_chany_bottom_out;
  wire [0:19] cby_1__1__1_chany_top_out;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__20_ccff_tail;
  wire [0:19] cby_1__1__20_chany_bottom_out;
  wire [0:19] cby_1__1__20_chany_top_out;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__21_ccff_tail;
  wire [0:19] cby_1__1__21_chany_bottom_out;
  wire [0:19] cby_1__1__21_chany_top_out;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__22_ccff_tail;
  wire [0:19] cby_1__1__22_chany_bottom_out;
  wire [0:19] cby_1__1__22_chany_top_out;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__23_ccff_tail;
  wire [0:19] cby_1__1__23_chany_bottom_out;
  wire [0:19] cby_1__1__23_chany_top_out;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__24_ccff_tail;
  wire [0:19] cby_1__1__24_chany_bottom_out;
  wire [0:19] cby_1__1__24_chany_top_out;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__25_ccff_tail;
  wire [0:19] cby_1__1__25_chany_bottom_out;
  wire [0:19] cby_1__1__25_chany_top_out;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__26_ccff_tail;
  wire [0:19] cby_1__1__26_chany_bottom_out;
  wire [0:19] cby_1__1__26_chany_top_out;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__27_ccff_tail;
  wire [0:19] cby_1__1__27_chany_bottom_out;
  wire [0:19] cby_1__1__27_chany_top_out;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__28_ccff_tail;
  wire [0:19] cby_1__1__28_chany_bottom_out;
  wire [0:19] cby_1__1__28_chany_top_out;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__29_ccff_tail;
  wire [0:19] cby_1__1__29_chany_bottom_out;
  wire [0:19] cby_1__1__29_chany_top_out;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__2_ccff_tail;
  wire [0:19] cby_1__1__2_chany_bottom_out;
  wire [0:19] cby_1__1__2_chany_top_out;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__30_ccff_tail;
  wire [0:19] cby_1__1__30_chany_bottom_out;
  wire [0:19] cby_1__1__30_chany_top_out;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__31_ccff_tail;
  wire [0:19] cby_1__1__31_chany_bottom_out;
  wire [0:19] cby_1__1__31_chany_top_out;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__32_ccff_tail;
  wire [0:19] cby_1__1__32_chany_bottom_out;
  wire [0:19] cby_1__1__32_chany_top_out;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__33_ccff_tail;
  wire [0:19] cby_1__1__33_chany_bottom_out;
  wire [0:19] cby_1__1__33_chany_top_out;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__34_ccff_tail;
  wire [0:19] cby_1__1__34_chany_bottom_out;
  wire [0:19] cby_1__1__34_chany_top_out;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__35_ccff_tail;
  wire [0:19] cby_1__1__35_chany_bottom_out;
  wire [0:19] cby_1__1__35_chany_top_out;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__36_ccff_tail;
  wire [0:19] cby_1__1__36_chany_bottom_out;
  wire [0:19] cby_1__1__36_chany_top_out;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__37_ccff_tail;
  wire [0:19] cby_1__1__37_chany_bottom_out;
  wire [0:19] cby_1__1__37_chany_top_out;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__38_ccff_tail;
  wire [0:19] cby_1__1__38_chany_bottom_out;
  wire [0:19] cby_1__1__38_chany_top_out;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__39_ccff_tail;
  wire [0:19] cby_1__1__39_chany_bottom_out;
  wire [0:19] cby_1__1__39_chany_top_out;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__3_ccff_tail;
  wire [0:19] cby_1__1__3_chany_bottom_out;
  wire [0:19] cby_1__1__3_chany_top_out;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__40_ccff_tail;
  wire [0:19] cby_1__1__40_chany_bottom_out;
  wire [0:19] cby_1__1__40_chany_top_out;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__41_ccff_tail;
  wire [0:19] cby_1__1__41_chany_bottom_out;
  wire [0:19] cby_1__1__41_chany_top_out;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__42_ccff_tail;
  wire [0:19] cby_1__1__42_chany_bottom_out;
  wire [0:19] cby_1__1__42_chany_top_out;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__43_ccff_tail;
  wire [0:19] cby_1__1__43_chany_bottom_out;
  wire [0:19] cby_1__1__43_chany_top_out;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__44_ccff_tail;
  wire [0:19] cby_1__1__44_chany_bottom_out;
  wire [0:19] cby_1__1__44_chany_top_out;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__45_ccff_tail;
  wire [0:19] cby_1__1__45_chany_bottom_out;
  wire [0:19] cby_1__1__45_chany_top_out;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__46_ccff_tail;
  wire [0:19] cby_1__1__46_chany_bottom_out;
  wire [0:19] cby_1__1__46_chany_top_out;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__47_ccff_tail;
  wire [0:19] cby_1__1__47_chany_bottom_out;
  wire [0:19] cby_1__1__47_chany_top_out;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__48_ccff_tail;
  wire [0:19] cby_1__1__48_chany_bottom_out;
  wire [0:19] cby_1__1__48_chany_top_out;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__49_ccff_tail;
  wire [0:19] cby_1__1__49_chany_bottom_out;
  wire [0:19] cby_1__1__49_chany_top_out;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__4_ccff_tail;
  wire [0:19] cby_1__1__4_chany_bottom_out;
  wire [0:19] cby_1__1__4_chany_top_out;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__50_ccff_tail;
  wire [0:19] cby_1__1__50_chany_bottom_out;
  wire [0:19] cby_1__1__50_chany_top_out;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__51_ccff_tail;
  wire [0:19] cby_1__1__51_chany_bottom_out;
  wire [0:19] cby_1__1__51_chany_top_out;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__52_ccff_tail;
  wire [0:19] cby_1__1__52_chany_bottom_out;
  wire [0:19] cby_1__1__52_chany_top_out;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__53_ccff_tail;
  wire [0:19] cby_1__1__53_chany_bottom_out;
  wire [0:19] cby_1__1__53_chany_top_out;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__54_ccff_tail;
  wire [0:19] cby_1__1__54_chany_bottom_out;
  wire [0:19] cby_1__1__54_chany_top_out;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__55_ccff_tail;
  wire [0:19] cby_1__1__55_chany_bottom_out;
  wire [0:19] cby_1__1__55_chany_top_out;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__56_ccff_tail;
  wire [0:19] cby_1__1__56_chany_bottom_out;
  wire [0:19] cby_1__1__56_chany_top_out;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__57_ccff_tail;
  wire [0:19] cby_1__1__57_chany_bottom_out;
  wire [0:19] cby_1__1__57_chany_top_out;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__58_ccff_tail;
  wire [0:19] cby_1__1__58_chany_bottom_out;
  wire [0:19] cby_1__1__58_chany_top_out;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__59_ccff_tail;
  wire [0:19] cby_1__1__59_chany_bottom_out;
  wire [0:19] cby_1__1__59_chany_top_out;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__5_ccff_tail;
  wire [0:19] cby_1__1__5_chany_bottom_out;
  wire [0:19] cby_1__1__5_chany_top_out;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__60_ccff_tail;
  wire [0:19] cby_1__1__60_chany_bottom_out;
  wire [0:19] cby_1__1__60_chany_top_out;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__61_ccff_tail;
  wire [0:19] cby_1__1__61_chany_bottom_out;
  wire [0:19] cby_1__1__61_chany_top_out;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__62_ccff_tail;
  wire [0:19] cby_1__1__62_chany_bottom_out;
  wire [0:19] cby_1__1__62_chany_top_out;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__63_ccff_tail;
  wire [0:19] cby_1__1__63_chany_bottom_out;
  wire [0:19] cby_1__1__63_chany_top_out;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__64_ccff_tail;
  wire [0:19] cby_1__1__64_chany_bottom_out;
  wire [0:19] cby_1__1__64_chany_top_out;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__65_ccff_tail;
  wire [0:19] cby_1__1__65_chany_bottom_out;
  wire [0:19] cby_1__1__65_chany_top_out;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__66_ccff_tail;
  wire [0:19] cby_1__1__66_chany_bottom_out;
  wire [0:19] cby_1__1__66_chany_top_out;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__67_ccff_tail;
  wire [0:19] cby_1__1__67_chany_bottom_out;
  wire [0:19] cby_1__1__67_chany_top_out;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__68_ccff_tail;
  wire [0:19] cby_1__1__68_chany_bottom_out;
  wire [0:19] cby_1__1__68_chany_top_out;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__69_ccff_tail;
  wire [0:19] cby_1__1__69_chany_bottom_out;
  wire [0:19] cby_1__1__69_chany_top_out;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__6_ccff_tail;
  wire [0:19] cby_1__1__6_chany_bottom_out;
  wire [0:19] cby_1__1__6_chany_top_out;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__70_ccff_tail;
  wire [0:19] cby_1__1__70_chany_bottom_out;
  wire [0:19] cby_1__1__70_chany_top_out;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__71_ccff_tail;
  wire [0:19] cby_1__1__71_chany_bottom_out;
  wire [0:19] cby_1__1__71_chany_top_out;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__72_ccff_tail;
  wire [0:19] cby_1__1__72_chany_bottom_out;
  wire [0:19] cby_1__1__72_chany_top_out;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__73_ccff_tail;
  wire [0:19] cby_1__1__73_chany_bottom_out;
  wire [0:19] cby_1__1__73_chany_top_out;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__74_ccff_tail;
  wire [0:19] cby_1__1__74_chany_bottom_out;
  wire [0:19] cby_1__1__74_chany_top_out;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__75_ccff_tail;
  wire [0:19] cby_1__1__75_chany_bottom_out;
  wire [0:19] cby_1__1__75_chany_top_out;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__76_ccff_tail;
  wire [0:19] cby_1__1__76_chany_bottom_out;
  wire [0:19] cby_1__1__76_chany_top_out;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__77_ccff_tail;
  wire [0:19] cby_1__1__77_chany_bottom_out;
  wire [0:19] cby_1__1__77_chany_top_out;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__78_ccff_tail;
  wire [0:19] cby_1__1__78_chany_bottom_out;
  wire [0:19] cby_1__1__78_chany_top_out;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__79_ccff_tail;
  wire [0:19] cby_1__1__79_chany_bottom_out;
  wire [0:19] cby_1__1__79_chany_top_out;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__7_ccff_tail;
  wire [0:19] cby_1__1__7_chany_bottom_out;
  wire [0:19] cby_1__1__7_chany_top_out;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__80_ccff_tail;
  wire [0:19] cby_1__1__80_chany_bottom_out;
  wire [0:19] cby_1__1__80_chany_top_out;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__81_ccff_tail;
  wire [0:19] cby_1__1__81_chany_bottom_out;
  wire [0:19] cby_1__1__81_chany_top_out;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__82_ccff_tail;
  wire [0:19] cby_1__1__82_chany_bottom_out;
  wire [0:19] cby_1__1__82_chany_top_out;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__83_ccff_tail;
  wire [0:19] cby_1__1__83_chany_bottom_out;
  wire [0:19] cby_1__1__83_chany_top_out;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__84_ccff_tail;
  wire [0:19] cby_1__1__84_chany_bottom_out;
  wire [0:19] cby_1__1__84_chany_top_out;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__85_ccff_tail;
  wire [0:19] cby_1__1__85_chany_bottom_out;
  wire [0:19] cby_1__1__85_chany_top_out;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__86_ccff_tail;
  wire [0:19] cby_1__1__86_chany_bottom_out;
  wire [0:19] cby_1__1__86_chany_top_out;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__87_ccff_tail;
  wire [0:19] cby_1__1__87_chany_bottom_out;
  wire [0:19] cby_1__1__87_chany_top_out;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__88_ccff_tail;
  wire [0:19] cby_1__1__88_chany_bottom_out;
  wire [0:19] cby_1__1__88_chany_top_out;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__89_ccff_tail;
  wire [0:19] cby_1__1__89_chany_bottom_out;
  wire [0:19] cby_1__1__89_chany_top_out;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__8_ccff_tail;
  wire [0:19] cby_1__1__8_chany_bottom_out;
  wire [0:19] cby_1__1__8_chany_top_out;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__90_ccff_tail;
  wire [0:19] cby_1__1__90_chany_bottom_out;
  wire [0:19] cby_1__1__90_chany_top_out;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__91_ccff_tail;
  wire [0:19] cby_1__1__91_chany_bottom_out;
  wire [0:19] cby_1__1__91_chany_top_out;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__92_ccff_tail;
  wire [0:19] cby_1__1__92_chany_bottom_out;
  wire [0:19] cby_1__1__92_chany_top_out;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__93_ccff_tail;
  wire [0:19] cby_1__1__93_chany_bottom_out;
  wire [0:19] cby_1__1__93_chany_top_out;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__94_ccff_tail;
  wire [0:19] cby_1__1__94_chany_bottom_out;
  wire [0:19] cby_1__1__94_chany_top_out;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__95_ccff_tail;
  wire [0:19] cby_1__1__95_chany_bottom_out;
  wire [0:19] cby_1__1__95_chany_top_out;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__96_ccff_tail;
  wire [0:19] cby_1__1__96_chany_bottom_out;
  wire [0:19] cby_1__1__96_chany_top_out;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__97_ccff_tail;
  wire [0:19] cby_1__1__97_chany_bottom_out;
  wire [0:19] cby_1__1__97_chany_top_out;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__98_ccff_tail;
  wire [0:19] cby_1__1__98_chany_bottom_out;
  wire [0:19] cby_1__1__98_chany_top_out;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__99_ccff_tail;
  wire [0:19] cby_1__1__99_chany_bottom_out;
  wire [0:19] cby_1__1__99_chany_top_out;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__9_ccff_tail;
  wire [0:19] cby_1__1__9_chany_bottom_out;
  wire [0:19] cby_1__1__9_chany_top_out;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:19] cby_1__3__0_chany_bottom_out;
  wire [0:19] cby_1__3__0_chany_top_out;
  wire [0:19] cby_1__3__10_chany_bottom_out;
  wire [0:19] cby_1__3__10_chany_top_out;
  wire [0:19] cby_1__3__11_chany_bottom_out;
  wire [0:19] cby_1__3__11_chany_top_out;
  wire [0:19] cby_1__3__1_chany_bottom_out;
  wire [0:19] cby_1__3__1_chany_top_out;
  wire [0:19] cby_1__3__2_chany_bottom_out;
  wire [0:19] cby_1__3__2_chany_top_out;
  wire [0:19] cby_1__3__3_chany_bottom_out;
  wire [0:19] cby_1__3__3_chany_top_out;
  wire [0:19] cby_1__3__4_chany_bottom_out;
  wire [0:19] cby_1__3__4_chany_top_out;
  wire [0:19] cby_1__3__5_chany_bottom_out;
  wire [0:19] cby_1__3__5_chany_top_out;
  wire [0:19] cby_1__3__6_chany_bottom_out;
  wire [0:19] cby_1__3__6_chany_top_out;
  wire [0:19] cby_1__3__7_chany_bottom_out;
  wire [0:19] cby_1__3__7_chany_top_out;
  wire [0:19] cby_1__3__8_chany_bottom_out;
  wire [0:19] cby_1__3__8_chany_top_out;
  wire [0:19] cby_1__3__9_chany_bottom_out;
  wire [0:19] cby_1__3__9_chany_top_out;
  wire [0:0] cby_2__3__0_ccff_tail;
  wire [0:19] cby_2__3__0_chany_bottom_out;
  wire [0:19] cby_2__3__0_chany_top_out;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__1_ccff_tail;
  wire [0:19] cby_2__3__1_chany_bottom_out;
  wire [0:19] cby_2__3__1_chany_top_out;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__2_ccff_tail;
  wire [0:19] cby_2__3__2_chany_bottom_out;
  wire [0:19] cby_2__3__2_chany_top_out;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__3_ccff_tail;
  wire [0:19] cby_2__3__3_chany_bottom_out;
  wire [0:19] cby_2__3__3_chany_top_out;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__4_ccff_tail;
  wire [0:19] cby_2__3__4_chany_bottom_out;
  wire [0:19] cby_2__3__4_chany_top_out;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__5_ccff_tail;
  wire [0:19] cby_2__3__5_chany_bottom_out;
  wire [0:19] cby_2__3__5_chany_top_out;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__6_ccff_tail;
  wire [0:19] cby_2__3__6_chany_bottom_out;
  wire [0:19] cby_2__3__6_chany_top_out;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__7_ccff_tail;
  wire [0:19] cby_2__3__7_chany_bottom_out;
  wire [0:19] cby_2__3__7_chany_top_out;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__8_ccff_tail;
  wire [0:19] cby_2__3__8_chany_bottom_out;
  wire [0:19] cby_2__3__8_chany_top_out;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__9_ccff_tail;
  wire [0:19] cby_2__3__9_chany_bottom_out;
  wire [0:19] cby_2__3__9_chany_top_out;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] direct_interc_0_out;
  wire [0:0] direct_interc_100_out;
  wire [0:0] direct_interc_101_out;
  wire [0:0] direct_interc_102_out;
  wire [0:0] direct_interc_103_out;
  wire [0:0] direct_interc_104_out;
  wire [0:0] direct_interc_105_out;
  wire [0:0] direct_interc_106_out;
  wire [0:0] direct_interc_107_out;
  wire [0:0] direct_interc_108_out;
  wire [0:0] direct_interc_109_out;
  wire [0:0] direct_interc_10_out;
  wire [0:0] direct_interc_110_out;
  wire [0:0] direct_interc_111_out;
  wire [0:0] direct_interc_112_out;
  wire [0:0] direct_interc_113_out;
  wire [0:0] direct_interc_114_out;
  wire [0:0] direct_interc_115_out;
  wire [0:0] direct_interc_116_out;
  wire [0:0] direct_interc_117_out;
  wire [0:0] direct_interc_118_out;
  wire [0:0] direct_interc_119_out;
  wire [0:0] direct_interc_11_out;
  wire [0:0] direct_interc_120_out;
  wire [0:0] direct_interc_121_out;
  wire [0:0] direct_interc_122_out;
  wire [0:0] direct_interc_123_out;
  wire [0:0] direct_interc_124_out;
  wire [0:0] direct_interc_125_out;
  wire [0:0] direct_interc_126_out;
  wire [0:0] direct_interc_127_out;
  wire [0:0] direct_interc_128_out;
  wire [0:0] direct_interc_129_out;
  wire [0:0] direct_interc_12_out;
  wire [0:0] direct_interc_130_out;
  wire [0:0] direct_interc_131_out;
  wire [0:0] direct_interc_132_out;
  wire [0:0] direct_interc_133_out;
  wire [0:0] direct_interc_134_out;
  wire [0:0] direct_interc_135_out;
  wire [0:0] direct_interc_136_out;
  wire [0:0] direct_interc_137_out;
  wire [0:0] direct_interc_138_out;
  wire [0:0] direct_interc_139_out;
  wire [0:0] direct_interc_13_out;
  wire [0:0] direct_interc_140_out;
  wire [0:0] direct_interc_141_out;
  wire [0:0] direct_interc_142_out;
  wire [0:0] direct_interc_143_out;
  wire [0:0] direct_interc_144_out;
  wire [0:0] direct_interc_145_out;
  wire [0:0] direct_interc_146_out;
  wire [0:0] direct_interc_147_out;
  wire [0:0] direct_interc_148_out;
  wire [0:0] direct_interc_149_out;
  wire [0:0] direct_interc_14_out;
  wire [0:0] direct_interc_150_out;
  wire [0:0] direct_interc_151_out;
  wire [0:0] direct_interc_152_out;
  wire [0:0] direct_interc_153_out;
  wire [0:0] direct_interc_154_out;
  wire [0:0] direct_interc_155_out;
  wire [0:0] direct_interc_156_out;
  wire [0:0] direct_interc_157_out;
  wire [0:0] direct_interc_158_out;
  wire [0:0] direct_interc_159_out;
  wire [0:0] direct_interc_15_out;
  wire [0:0] direct_interc_160_out;
  wire [0:0] direct_interc_161_out;
  wire [0:0] direct_interc_162_out;
  wire [0:0] direct_interc_163_out;
  wire [0:0] direct_interc_164_out;
  wire [0:0] direct_interc_165_out;
  wire [0:0] direct_interc_166_out;
  wire [0:0] direct_interc_167_out;
  wire [0:0] direct_interc_168_out;
  wire [0:0] direct_interc_169_out;
  wire [0:0] direct_interc_16_out;
  wire [0:0] direct_interc_170_out;
  wire [0:0] direct_interc_171_out;
  wire [0:0] direct_interc_172_out;
  wire [0:0] direct_interc_173_out;
  wire [0:0] direct_interc_174_out;
  wire [0:0] direct_interc_175_out;
  wire [0:0] direct_interc_176_out;
  wire [0:0] direct_interc_177_out;
  wire [0:0] direct_interc_178_out;
  wire [0:0] direct_interc_17_out;
  wire [0:0] direct_interc_18_out;
  wire [0:0] direct_interc_19_out;
  wire [0:0] direct_interc_1_out;
  wire [0:0] direct_interc_20_out;
  wire [0:0] direct_interc_21_out;
  wire [0:0] direct_interc_22_out;
  wire [0:0] direct_interc_23_out;
  wire [0:0] direct_interc_24_out;
  wire [0:0] direct_interc_25_out;
  wire [0:0] direct_interc_26_out;
  wire [0:0] direct_interc_27_out;
  wire [0:0] direct_interc_28_out;
  wire [0:0] direct_interc_29_out;
  wire [0:0] direct_interc_2_out;
  wire [0:0] direct_interc_30_out;
  wire [0:0] direct_interc_31_out;
  wire [0:0] direct_interc_32_out;
  wire [0:0] direct_interc_33_out;
  wire [0:0] direct_interc_34_out;
  wire [0:0] direct_interc_35_out;
  wire [0:0] direct_interc_36_out;
  wire [0:0] direct_interc_37_out;
  wire [0:0] direct_interc_38_out;
  wire [0:0] direct_interc_39_out;
  wire [0:0] direct_interc_3_out;
  wire [0:0] direct_interc_40_out;
  wire [0:0] direct_interc_41_out;
  wire [0:0] direct_interc_42_out;
  wire [0:0] direct_interc_43_out;
  wire [0:0] direct_interc_44_out;
  wire [0:0] direct_interc_45_out;
  wire [0:0] direct_interc_46_out;
  wire [0:0] direct_interc_47_out;
  wire [0:0] direct_interc_48_out;
  wire [0:0] direct_interc_49_out;
  wire [0:0] direct_interc_4_out;
  wire [0:0] direct_interc_50_out;
  wire [0:0] direct_interc_51_out;
  wire [0:0] direct_interc_52_out;
  wire [0:0] direct_interc_53_out;
  wire [0:0] direct_interc_54_out;
  wire [0:0] direct_interc_55_out;
  wire [0:0] direct_interc_56_out;
  wire [0:0] direct_interc_57_out;
  wire [0:0] direct_interc_58_out;
  wire [0:0] direct_interc_59_out;
  wire [0:0] direct_interc_5_out;
  wire [0:0] direct_interc_60_out;
  wire [0:0] direct_interc_61_out;
  wire [0:0] direct_interc_62_out;
  wire [0:0] direct_interc_63_out;
  wire [0:0] direct_interc_64_out;
  wire [0:0] direct_interc_65_out;
  wire [0:0] direct_interc_66_out;
  wire [0:0] direct_interc_67_out;
  wire [0:0] direct_interc_68_out;
  wire [0:0] direct_interc_69_out;
  wire [0:0] direct_interc_6_out;
  wire [0:0] direct_interc_70_out;
  wire [0:0] direct_interc_71_out;
  wire [0:0] direct_interc_72_out;
  wire [0:0] direct_interc_73_out;
  wire [0:0] direct_interc_74_out;
  wire [0:0] direct_interc_75_out;
  wire [0:0] direct_interc_76_out;
  wire [0:0] direct_interc_77_out;
  wire [0:0] direct_interc_78_out;
  wire [0:0] direct_interc_79_out;
  wire [0:0] direct_interc_7_out;
  wire [0:0] direct_interc_80_out;
  wire [0:0] direct_interc_81_out;
  wire [0:0] direct_interc_82_out;
  wire [0:0] direct_interc_83_out;
  wire [0:0] direct_interc_84_out;
  wire [0:0] direct_interc_85_out;
  wire [0:0] direct_interc_86_out;
  wire [0:0] direct_interc_87_out;
  wire [0:0] direct_interc_88_out;
  wire [0:0] direct_interc_89_out;
  wire [0:0] direct_interc_8_out;
  wire [0:0] direct_interc_90_out;
  wire [0:0] direct_interc_91_out;
  wire [0:0] direct_interc_92_out;
  wire [0:0] direct_interc_93_out;
  wire [0:0] direct_interc_94_out;
  wire [0:0] direct_interc_95_out;
  wire [0:0] direct_interc_96_out;
  wire [0:0] direct_interc_97_out;
  wire [0:0] direct_interc_98_out;
  wire [0:0] direct_interc_99_out;
  wire [0:0] direct_interc_9_out;
  wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_0_ccff_tail;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_100_ccff_tail;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_101_ccff_tail;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_102_ccff_tail;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_103_ccff_tail;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_104_ccff_tail;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_105_ccff_tail;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_106_ccff_tail;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_107_ccff_tail;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_108_ccff_tail;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_109_ccff_tail;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10_ccff_tail;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_110_ccff_tail;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_111_ccff_tail;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_112_ccff_tail;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_113_ccff_tail;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_114_ccff_tail;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_115_ccff_tail;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_116_ccff_tail;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_117_ccff_tail;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_118_ccff_tail;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_119_ccff_tail;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11_ccff_tail;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_12_ccff_tail;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_13_ccff_tail;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_14_ccff_tail;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_15_ccff_tail;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_16_ccff_tail;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_17_ccff_tail;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_18_ccff_tail;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_19_ccff_tail;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1_ccff_tail;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_20_ccff_tail;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_21_ccff_tail;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_22_ccff_tail;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_23_ccff_tail;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_24_ccff_tail;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_25_ccff_tail;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_26_ccff_tail;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_27_ccff_tail;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_28_ccff_tail;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_29_ccff_tail;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_2__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_2_ccff_tail;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_30_ccff_tail;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_31_ccff_tail;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_32_ccff_tail;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_33_ccff_tail;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_34_ccff_tail;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_35_ccff_tail;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_36_ccff_tail;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_37_ccff_tail;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_38_ccff_tail;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_39_ccff_tail;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3_ccff_tail;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_40_ccff_tail;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_41_ccff_tail;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_42_ccff_tail;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_43_ccff_tail;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_44_ccff_tail;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_45_ccff_tail;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_46_ccff_tail;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_47_ccff_tail;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_48_ccff_tail;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_49_ccff_tail;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4_ccff_tail;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_50_ccff_tail;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_51_ccff_tail;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_52_ccff_tail;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_53_ccff_tail;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_54_ccff_tail;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_55_ccff_tail;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_56_ccff_tail;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_57_ccff_tail;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_58_ccff_tail;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_59_ccff_tail;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5_ccff_tail;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_60_ccff_tail;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_61_ccff_tail;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_62_ccff_tail;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_63_ccff_tail;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_64_ccff_tail;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_65_ccff_tail;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_66_ccff_tail;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_67_ccff_tail;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_68_ccff_tail;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_69_ccff_tail;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6_ccff_tail;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_70_ccff_tail;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_71_ccff_tail;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_72_ccff_tail;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_73_ccff_tail;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_74_ccff_tail;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_75_ccff_tail;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_76_ccff_tail;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_77_ccff_tail;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_78_ccff_tail;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_79_ccff_tail;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7_ccff_tail;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_80_ccff_tail;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_81_ccff_tail;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_82_ccff_tail;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_83_ccff_tail;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_84_ccff_tail;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_85_ccff_tail;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_86_ccff_tail;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_87_ccff_tail;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_88_ccff_tail;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_89_ccff_tail;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_8__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_8_ccff_tail;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_90_ccff_tail;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_91_ccff_tail;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_92_ccff_tail;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_93_ccff_tail;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_94_ccff_tail;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_95_ccff_tail;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_96_ccff_tail;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_97_ccff_tail;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_98_ccff_tail;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_99_ccff_tail;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9_ccff_tail;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_0_ccff_tail;
  wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_10_ccff_tail;
  wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_11_ccff_tail;
  wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_1_ccff_tail;
  wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_2_ccff_tail;
  wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_3_ccff_tail;
  wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_4_ccff_tail;
  wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_5_ccff_tail;
  wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_6_ccff_tail;
  wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_7_ccff_tail;
  wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_8_ccff_tail;
  wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_9_ccff_tail;
  wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_0_ccff_tail;
  wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_10_ccff_tail;
  wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_11_ccff_tail;
  wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_1_ccff_tail;
  wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_2_ccff_tail;
  wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_3_ccff_tail;
  wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_4_ccff_tail;
  wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_5_ccff_tail;
  wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_6_ccff_tail;
  wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_7_ccff_tail;
  wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_8_ccff_tail;
  wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_9_ccff_tail;
  wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_0_ccff_tail;
  wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_10_ccff_tail;
  wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_11_ccff_tail;
  wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_1_ccff_tail;
  wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_2_ccff_tail;
  wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_3_ccff_tail;
  wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_4_ccff_tail;
  wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_5_ccff_tail;
  wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_6_ccff_tail;
  wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_7_ccff_tail;
  wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_8_ccff_tail;
  wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_9_ccff_tail;
  wire [0:0] grid_mult_18_0_ccff_tail;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_10_ccff_tail;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_11_ccff_tail;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_1_ccff_tail;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_2_ccff_tail;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_3_ccff_tail;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_4_ccff_tail;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_5_ccff_tail;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_6_ccff_tail;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_7_ccff_tail;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_8_ccff_tail;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_9_ccff_tail;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] sb_0__0__0_ccff_tail;
  wire [0:19] sb_0__0__0_chanx_right_out;
  wire [0:19] sb_0__0__0_chany_top_out;
  wire [0:0] sb_0__12__0_ccff_tail;
  wire [0:19] sb_0__12__0_chanx_right_out;
  wire [0:19] sb_0__12__0_chany_bottom_out;
  wire [0:0] sb_0__1__0_ccff_tail;
  wire [0:19] sb_0__1__0_chanx_right_out;
  wire [0:19] sb_0__1__0_chany_bottom_out;
  wire [0:19] sb_0__1__0_chany_top_out;
  wire [0:0] sb_0__1__1_ccff_tail;
  wire [0:19] sb_0__1__1_chanx_right_out;
  wire [0:19] sb_0__1__1_chany_bottom_out;
  wire [0:19] sb_0__1__1_chany_top_out;
  wire [0:0] sb_0__1__2_ccff_tail;
  wire [0:19] sb_0__1__2_chanx_right_out;
  wire [0:19] sb_0__1__2_chany_bottom_out;
  wire [0:19] sb_0__1__2_chany_top_out;
  wire [0:0] sb_0__1__3_ccff_tail;
  wire [0:19] sb_0__1__3_chanx_right_out;
  wire [0:19] sb_0__1__3_chany_bottom_out;
  wire [0:19] sb_0__1__3_chany_top_out;
  wire [0:0] sb_0__1__4_ccff_tail;
  wire [0:19] sb_0__1__4_chanx_right_out;
  wire [0:19] sb_0__1__4_chany_bottom_out;
  wire [0:19] sb_0__1__4_chany_top_out;
  wire [0:0] sb_0__1__5_ccff_tail;
  wire [0:19] sb_0__1__5_chanx_right_out;
  wire [0:19] sb_0__1__5_chany_bottom_out;
  wire [0:19] sb_0__1__5_chany_top_out;
  wire [0:0] sb_0__1__6_ccff_tail;
  wire [0:19] sb_0__1__6_chanx_right_out;
  wire [0:19] sb_0__1__6_chany_bottom_out;
  wire [0:19] sb_0__1__6_chany_top_out;
  wire [0:0] sb_0__1__7_ccff_tail;
  wire [0:19] sb_0__1__7_chanx_right_out;
  wire [0:19] sb_0__1__7_chany_bottom_out;
  wire [0:19] sb_0__1__7_chany_top_out;
  wire [0:0] sb_0__1__8_ccff_tail;
  wire [0:19] sb_0__1__8_chanx_right_out;
  wire [0:19] sb_0__1__8_chany_bottom_out;
  wire [0:19] sb_0__1__8_chany_top_out;
  wire [0:0] sb_0__3__0_ccff_tail;
  wire [0:19] sb_0__3__0_chanx_right_out;
  wire [0:19] sb_0__3__0_chany_bottom_out;
  wire [0:19] sb_0__3__0_chany_top_out;
  wire [0:0] sb_0__3__1_ccff_tail;
  wire [0:19] sb_0__3__1_chanx_right_out;
  wire [0:19] sb_0__3__1_chany_bottom_out;
  wire [0:19] sb_0__3__1_chany_top_out;
  wire [0:19] sb_12__0__0_chanx_left_out;
  wire [0:19] sb_12__0__0_chany_top_out;
  wire [0:0] sb_12__12__0_ccff_tail;
  wire [0:19] sb_12__12__0_chanx_left_out;
  wire [0:19] sb_12__12__0_chany_bottom_out;
  wire [0:19] sb_12__1__0_chanx_left_out;
  wire [0:19] sb_12__1__0_chany_bottom_out;
  wire [0:19] sb_12__1__0_chany_top_out;
  wire [0:19] sb_12__1__1_chanx_left_out;
  wire [0:19] sb_12__1__1_chany_bottom_out;
  wire [0:19] sb_12__1__1_chany_top_out;
  wire [0:19] sb_12__1__2_chanx_left_out;
  wire [0:19] sb_12__1__2_chany_bottom_out;
  wire [0:19] sb_12__1__2_chany_top_out;
  wire [0:19] sb_12__1__3_chanx_left_out;
  wire [0:19] sb_12__1__3_chany_bottom_out;
  wire [0:19] sb_12__1__3_chany_top_out;
  wire [0:19] sb_12__1__4_chanx_left_out;
  wire [0:19] sb_12__1__4_chany_bottom_out;
  wire [0:19] sb_12__1__4_chany_top_out;
  wire [0:19] sb_12__1__5_chanx_left_out;
  wire [0:19] sb_12__1__5_chany_bottom_out;
  wire [0:19] sb_12__1__5_chany_top_out;
  wire [0:19] sb_12__1__6_chanx_left_out;
  wire [0:19] sb_12__1__6_chany_bottom_out;
  wire [0:19] sb_12__1__6_chany_top_out;
  wire [0:19] sb_12__2__0_chanx_left_out;
  wire [0:19] sb_12__2__0_chany_bottom_out;
  wire [0:19] sb_12__2__0_chany_top_out;
  wire [0:19] sb_12__2__1_chanx_left_out;
  wire [0:19] sb_12__2__1_chany_bottom_out;
  wire [0:19] sb_12__2__1_chany_top_out;
  wire [0:19] sb_12__3__0_chanx_left_out;
  wire [0:19] sb_12__3__0_chany_bottom_out;
  wire [0:19] sb_12__3__0_chany_top_out;
  wire [0:19] sb_12__3__1_chanx_left_out;
  wire [0:19] sb_12__3__1_chany_bottom_out;
  wire [0:19] sb_12__3__1_chany_top_out;
  wire [0:0] sb_1__0__0_ccff_tail;
  wire [0:19] sb_1__0__0_chanx_left_out;
  wire [0:19] sb_1__0__0_chanx_right_out;
  wire [0:19] sb_1__0__0_chany_top_out;
  wire [0:0] sb_1__0__10_ccff_tail;
  wire [0:19] sb_1__0__10_chanx_left_out;
  wire [0:19] sb_1__0__10_chanx_right_out;
  wire [0:19] sb_1__0__10_chany_top_out;
  wire [0:0] sb_1__0__1_ccff_tail;
  wire [0:19] sb_1__0__1_chanx_left_out;
  wire [0:19] sb_1__0__1_chanx_right_out;
  wire [0:19] sb_1__0__1_chany_top_out;
  wire [0:0] sb_1__0__2_ccff_tail;
  wire [0:19] sb_1__0__2_chanx_left_out;
  wire [0:19] sb_1__0__2_chanx_right_out;
  wire [0:19] sb_1__0__2_chany_top_out;
  wire [0:0] sb_1__0__3_ccff_tail;
  wire [0:19] sb_1__0__3_chanx_left_out;
  wire [0:19] sb_1__0__3_chanx_right_out;
  wire [0:19] sb_1__0__3_chany_top_out;
  wire [0:0] sb_1__0__4_ccff_tail;
  wire [0:19] sb_1__0__4_chanx_left_out;
  wire [0:19] sb_1__0__4_chanx_right_out;
  wire [0:19] sb_1__0__4_chany_top_out;
  wire [0:0] sb_1__0__5_ccff_tail;
  wire [0:19] sb_1__0__5_chanx_left_out;
  wire [0:19] sb_1__0__5_chanx_right_out;
  wire [0:19] sb_1__0__5_chany_top_out;
  wire [0:0] sb_1__0__6_ccff_tail;
  wire [0:19] sb_1__0__6_chanx_left_out;
  wire [0:19] sb_1__0__6_chanx_right_out;
  wire [0:19] sb_1__0__6_chany_top_out;
  wire [0:0] sb_1__0__7_ccff_tail;
  wire [0:19] sb_1__0__7_chanx_left_out;
  wire [0:19] sb_1__0__7_chanx_right_out;
  wire [0:19] sb_1__0__7_chany_top_out;
  wire [0:0] sb_1__0__8_ccff_tail;
  wire [0:19] sb_1__0__8_chanx_left_out;
  wire [0:19] sb_1__0__8_chanx_right_out;
  wire [0:19] sb_1__0__8_chany_top_out;
  wire [0:0] sb_1__0__9_ccff_tail;
  wire [0:19] sb_1__0__9_chanx_left_out;
  wire [0:19] sb_1__0__9_chanx_right_out;
  wire [0:19] sb_1__0__9_chany_top_out;
  wire [0:0] sb_1__12__0_ccff_tail;
  wire [0:19] sb_1__12__0_chanx_left_out;
  wire [0:19] sb_1__12__0_chanx_right_out;
  wire [0:19] sb_1__12__0_chany_bottom_out;
  wire [0:0] sb_1__12__10_ccff_tail;
  wire [0:19] sb_1__12__10_chanx_left_out;
  wire [0:19] sb_1__12__10_chanx_right_out;
  wire [0:19] sb_1__12__10_chany_bottom_out;
  wire [0:0] sb_1__12__1_ccff_tail;
  wire [0:19] sb_1__12__1_chanx_left_out;
  wire [0:19] sb_1__12__1_chanx_right_out;
  wire [0:19] sb_1__12__1_chany_bottom_out;
  wire [0:0] sb_1__12__2_ccff_tail;
  wire [0:19] sb_1__12__2_chanx_left_out;
  wire [0:19] sb_1__12__2_chanx_right_out;
  wire [0:19] sb_1__12__2_chany_bottom_out;
  wire [0:0] sb_1__12__3_ccff_tail;
  wire [0:19] sb_1__12__3_chanx_left_out;
  wire [0:19] sb_1__12__3_chanx_right_out;
  wire [0:19] sb_1__12__3_chany_bottom_out;
  wire [0:0] sb_1__12__4_ccff_tail;
  wire [0:19] sb_1__12__4_chanx_left_out;
  wire [0:19] sb_1__12__4_chanx_right_out;
  wire [0:19] sb_1__12__4_chany_bottom_out;
  wire [0:0] sb_1__12__5_ccff_tail;
  wire [0:19] sb_1__12__5_chanx_left_out;
  wire [0:19] sb_1__12__5_chanx_right_out;
  wire [0:19] sb_1__12__5_chany_bottom_out;
  wire [0:0] sb_1__12__6_ccff_tail;
  wire [0:19] sb_1__12__6_chanx_left_out;
  wire [0:19] sb_1__12__6_chanx_right_out;
  wire [0:19] sb_1__12__6_chany_bottom_out;
  wire [0:0] sb_1__12__7_ccff_tail;
  wire [0:19] sb_1__12__7_chanx_left_out;
  wire [0:19] sb_1__12__7_chanx_right_out;
  wire [0:19] sb_1__12__7_chany_bottom_out;
  wire [0:0] sb_1__12__8_ccff_tail;
  wire [0:19] sb_1__12__8_chanx_left_out;
  wire [0:19] sb_1__12__8_chanx_right_out;
  wire [0:19] sb_1__12__8_chany_bottom_out;
  wire [0:0] sb_1__12__9_ccff_tail;
  wire [0:19] sb_1__12__9_chanx_left_out;
  wire [0:19] sb_1__12__9_chanx_right_out;
  wire [0:19] sb_1__12__9_chany_bottom_out;
  wire [0:0] sb_1__1__0_ccff_tail;
  wire [0:19] sb_1__1__0_chanx_left_out;
  wire [0:19] sb_1__1__0_chanx_right_out;
  wire [0:19] sb_1__1__0_chany_bottom_out;
  wire [0:19] sb_1__1__0_chany_top_out;
  wire [0:0] sb_1__1__10_ccff_tail;
  wire [0:19] sb_1__1__10_chanx_left_out;
  wire [0:19] sb_1__1__10_chanx_right_out;
  wire [0:19] sb_1__1__10_chany_bottom_out;
  wire [0:19] sb_1__1__10_chany_top_out;
  wire [0:0] sb_1__1__11_ccff_tail;
  wire [0:19] sb_1__1__11_chanx_left_out;
  wire [0:19] sb_1__1__11_chanx_right_out;
  wire [0:19] sb_1__1__11_chany_bottom_out;
  wire [0:19] sb_1__1__11_chany_top_out;
  wire [0:0] sb_1__1__12_ccff_tail;
  wire [0:19] sb_1__1__12_chanx_left_out;
  wire [0:19] sb_1__1__12_chanx_right_out;
  wire [0:19] sb_1__1__12_chany_bottom_out;
  wire [0:19] sb_1__1__12_chany_top_out;
  wire [0:0] sb_1__1__13_ccff_tail;
  wire [0:19] sb_1__1__13_chanx_left_out;
  wire [0:19] sb_1__1__13_chanx_right_out;
  wire [0:19] sb_1__1__13_chany_bottom_out;
  wire [0:19] sb_1__1__13_chany_top_out;
  wire [0:0] sb_1__1__14_ccff_tail;
  wire [0:19] sb_1__1__14_chanx_left_out;
  wire [0:19] sb_1__1__14_chanx_right_out;
  wire [0:19] sb_1__1__14_chany_bottom_out;
  wire [0:19] sb_1__1__14_chany_top_out;
  wire [0:0] sb_1__1__15_ccff_tail;
  wire [0:19] sb_1__1__15_chanx_left_out;
  wire [0:19] sb_1__1__15_chanx_right_out;
  wire [0:19] sb_1__1__15_chany_bottom_out;
  wire [0:19] sb_1__1__15_chany_top_out;
  wire [0:0] sb_1__1__16_ccff_tail;
  wire [0:19] sb_1__1__16_chanx_left_out;
  wire [0:19] sb_1__1__16_chanx_right_out;
  wire [0:19] sb_1__1__16_chany_bottom_out;
  wire [0:19] sb_1__1__16_chany_top_out;
  wire [0:0] sb_1__1__17_ccff_tail;
  wire [0:19] sb_1__1__17_chanx_left_out;
  wire [0:19] sb_1__1__17_chanx_right_out;
  wire [0:19] sb_1__1__17_chany_bottom_out;
  wire [0:19] sb_1__1__17_chany_top_out;
  wire [0:0] sb_1__1__18_ccff_tail;
  wire [0:19] sb_1__1__18_chanx_left_out;
  wire [0:19] sb_1__1__18_chanx_right_out;
  wire [0:19] sb_1__1__18_chany_bottom_out;
  wire [0:19] sb_1__1__18_chany_top_out;
  wire [0:0] sb_1__1__19_ccff_tail;
  wire [0:19] sb_1__1__19_chanx_left_out;
  wire [0:19] sb_1__1__19_chanx_right_out;
  wire [0:19] sb_1__1__19_chany_bottom_out;
  wire [0:19] sb_1__1__19_chany_top_out;
  wire [0:0] sb_1__1__1_ccff_tail;
  wire [0:19] sb_1__1__1_chanx_left_out;
  wire [0:19] sb_1__1__1_chanx_right_out;
  wire [0:19] sb_1__1__1_chany_bottom_out;
  wire [0:19] sb_1__1__1_chany_top_out;
  wire [0:0] sb_1__1__20_ccff_tail;
  wire [0:19] sb_1__1__20_chanx_left_out;
  wire [0:19] sb_1__1__20_chanx_right_out;
  wire [0:19] sb_1__1__20_chany_bottom_out;
  wire [0:19] sb_1__1__20_chany_top_out;
  wire [0:0] sb_1__1__21_ccff_tail;
  wire [0:19] sb_1__1__21_chanx_left_out;
  wire [0:19] sb_1__1__21_chanx_right_out;
  wire [0:19] sb_1__1__21_chany_bottom_out;
  wire [0:19] sb_1__1__21_chany_top_out;
  wire [0:0] sb_1__1__22_ccff_tail;
  wire [0:19] sb_1__1__22_chanx_left_out;
  wire [0:19] sb_1__1__22_chanx_right_out;
  wire [0:19] sb_1__1__22_chany_bottom_out;
  wire [0:19] sb_1__1__22_chany_top_out;
  wire [0:0] sb_1__1__23_ccff_tail;
  wire [0:19] sb_1__1__23_chanx_left_out;
  wire [0:19] sb_1__1__23_chanx_right_out;
  wire [0:19] sb_1__1__23_chany_bottom_out;
  wire [0:19] sb_1__1__23_chany_top_out;
  wire [0:0] sb_1__1__24_ccff_tail;
  wire [0:19] sb_1__1__24_chanx_left_out;
  wire [0:19] sb_1__1__24_chanx_right_out;
  wire [0:19] sb_1__1__24_chany_bottom_out;
  wire [0:19] sb_1__1__24_chany_top_out;
  wire [0:0] sb_1__1__25_ccff_tail;
  wire [0:19] sb_1__1__25_chanx_left_out;
  wire [0:19] sb_1__1__25_chanx_right_out;
  wire [0:19] sb_1__1__25_chany_bottom_out;
  wire [0:19] sb_1__1__25_chany_top_out;
  wire [0:0] sb_1__1__26_ccff_tail;
  wire [0:19] sb_1__1__26_chanx_left_out;
  wire [0:19] sb_1__1__26_chanx_right_out;
  wire [0:19] sb_1__1__26_chany_bottom_out;
  wire [0:19] sb_1__1__26_chany_top_out;
  wire [0:0] sb_1__1__27_ccff_tail;
  wire [0:19] sb_1__1__27_chanx_left_out;
  wire [0:19] sb_1__1__27_chanx_right_out;
  wire [0:19] sb_1__1__27_chany_bottom_out;
  wire [0:19] sb_1__1__27_chany_top_out;
  wire [0:0] sb_1__1__28_ccff_tail;
  wire [0:19] sb_1__1__28_chanx_left_out;
  wire [0:19] sb_1__1__28_chanx_right_out;
  wire [0:19] sb_1__1__28_chany_bottom_out;
  wire [0:19] sb_1__1__28_chany_top_out;
  wire [0:0] sb_1__1__29_ccff_tail;
  wire [0:19] sb_1__1__29_chanx_left_out;
  wire [0:19] sb_1__1__29_chanx_right_out;
  wire [0:19] sb_1__1__29_chany_bottom_out;
  wire [0:19] sb_1__1__29_chany_top_out;
  wire [0:0] sb_1__1__2_ccff_tail;
  wire [0:19] sb_1__1__2_chanx_left_out;
  wire [0:19] sb_1__1__2_chanx_right_out;
  wire [0:19] sb_1__1__2_chany_bottom_out;
  wire [0:19] sb_1__1__2_chany_top_out;
  wire [0:0] sb_1__1__30_ccff_tail;
  wire [0:19] sb_1__1__30_chanx_left_out;
  wire [0:19] sb_1__1__30_chanx_right_out;
  wire [0:19] sb_1__1__30_chany_bottom_out;
  wire [0:19] sb_1__1__30_chany_top_out;
  wire [0:0] sb_1__1__31_ccff_tail;
  wire [0:19] sb_1__1__31_chanx_left_out;
  wire [0:19] sb_1__1__31_chanx_right_out;
  wire [0:19] sb_1__1__31_chany_bottom_out;
  wire [0:19] sb_1__1__31_chany_top_out;
  wire [0:0] sb_1__1__32_ccff_tail;
  wire [0:19] sb_1__1__32_chanx_left_out;
  wire [0:19] sb_1__1__32_chanx_right_out;
  wire [0:19] sb_1__1__32_chany_bottom_out;
  wire [0:19] sb_1__1__32_chany_top_out;
  wire [0:0] sb_1__1__33_ccff_tail;
  wire [0:19] sb_1__1__33_chanx_left_out;
  wire [0:19] sb_1__1__33_chanx_right_out;
  wire [0:19] sb_1__1__33_chany_bottom_out;
  wire [0:19] sb_1__1__33_chany_top_out;
  wire [0:0] sb_1__1__34_ccff_tail;
  wire [0:19] sb_1__1__34_chanx_left_out;
  wire [0:19] sb_1__1__34_chanx_right_out;
  wire [0:19] sb_1__1__34_chany_bottom_out;
  wire [0:19] sb_1__1__34_chany_top_out;
  wire [0:0] sb_1__1__35_ccff_tail;
  wire [0:19] sb_1__1__35_chanx_left_out;
  wire [0:19] sb_1__1__35_chanx_right_out;
  wire [0:19] sb_1__1__35_chany_bottom_out;
  wire [0:19] sb_1__1__35_chany_top_out;
  wire [0:0] sb_1__1__36_ccff_tail;
  wire [0:19] sb_1__1__36_chanx_left_out;
  wire [0:19] sb_1__1__36_chanx_right_out;
  wire [0:19] sb_1__1__36_chany_bottom_out;
  wire [0:19] sb_1__1__36_chany_top_out;
  wire [0:0] sb_1__1__37_ccff_tail;
  wire [0:19] sb_1__1__37_chanx_left_out;
  wire [0:19] sb_1__1__37_chanx_right_out;
  wire [0:19] sb_1__1__37_chany_bottom_out;
  wire [0:19] sb_1__1__37_chany_top_out;
  wire [0:0] sb_1__1__38_ccff_tail;
  wire [0:19] sb_1__1__38_chanx_left_out;
  wire [0:19] sb_1__1__38_chanx_right_out;
  wire [0:19] sb_1__1__38_chany_bottom_out;
  wire [0:19] sb_1__1__38_chany_top_out;
  wire [0:0] sb_1__1__39_ccff_tail;
  wire [0:19] sb_1__1__39_chanx_left_out;
  wire [0:19] sb_1__1__39_chanx_right_out;
  wire [0:19] sb_1__1__39_chany_bottom_out;
  wire [0:19] sb_1__1__39_chany_top_out;
  wire [0:0] sb_1__1__3_ccff_tail;
  wire [0:19] sb_1__1__3_chanx_left_out;
  wire [0:19] sb_1__1__3_chanx_right_out;
  wire [0:19] sb_1__1__3_chany_bottom_out;
  wire [0:19] sb_1__1__3_chany_top_out;
  wire [0:0] sb_1__1__40_ccff_tail;
  wire [0:19] sb_1__1__40_chanx_left_out;
  wire [0:19] sb_1__1__40_chanx_right_out;
  wire [0:19] sb_1__1__40_chany_bottom_out;
  wire [0:19] sb_1__1__40_chany_top_out;
  wire [0:0] sb_1__1__41_ccff_tail;
  wire [0:19] sb_1__1__41_chanx_left_out;
  wire [0:19] sb_1__1__41_chanx_right_out;
  wire [0:19] sb_1__1__41_chany_bottom_out;
  wire [0:19] sb_1__1__41_chany_top_out;
  wire [0:0] sb_1__1__42_ccff_tail;
  wire [0:19] sb_1__1__42_chanx_left_out;
  wire [0:19] sb_1__1__42_chanx_right_out;
  wire [0:19] sb_1__1__42_chany_bottom_out;
  wire [0:19] sb_1__1__42_chany_top_out;
  wire [0:0] sb_1__1__43_ccff_tail;
  wire [0:19] sb_1__1__43_chanx_left_out;
  wire [0:19] sb_1__1__43_chanx_right_out;
  wire [0:19] sb_1__1__43_chany_bottom_out;
  wire [0:19] sb_1__1__43_chany_top_out;
  wire [0:0] sb_1__1__44_ccff_tail;
  wire [0:19] sb_1__1__44_chanx_left_out;
  wire [0:19] sb_1__1__44_chanx_right_out;
  wire [0:19] sb_1__1__44_chany_bottom_out;
  wire [0:19] sb_1__1__44_chany_top_out;
  wire [0:0] sb_1__1__45_ccff_tail;
  wire [0:19] sb_1__1__45_chanx_left_out;
  wire [0:19] sb_1__1__45_chanx_right_out;
  wire [0:19] sb_1__1__45_chany_bottom_out;
  wire [0:19] sb_1__1__45_chany_top_out;
  wire [0:0] sb_1__1__46_ccff_tail;
  wire [0:19] sb_1__1__46_chanx_left_out;
  wire [0:19] sb_1__1__46_chanx_right_out;
  wire [0:19] sb_1__1__46_chany_bottom_out;
  wire [0:19] sb_1__1__46_chany_top_out;
  wire [0:0] sb_1__1__47_ccff_tail;
  wire [0:19] sb_1__1__47_chanx_left_out;
  wire [0:19] sb_1__1__47_chanx_right_out;
  wire [0:19] sb_1__1__47_chany_bottom_out;
  wire [0:19] sb_1__1__47_chany_top_out;
  wire [0:0] sb_1__1__48_ccff_tail;
  wire [0:19] sb_1__1__48_chanx_left_out;
  wire [0:19] sb_1__1__48_chanx_right_out;
  wire [0:19] sb_1__1__48_chany_bottom_out;
  wire [0:19] sb_1__1__48_chany_top_out;
  wire [0:0] sb_1__1__49_ccff_tail;
  wire [0:19] sb_1__1__49_chanx_left_out;
  wire [0:19] sb_1__1__49_chanx_right_out;
  wire [0:19] sb_1__1__49_chany_bottom_out;
  wire [0:19] sb_1__1__49_chany_top_out;
  wire [0:0] sb_1__1__4_ccff_tail;
  wire [0:19] sb_1__1__4_chanx_left_out;
  wire [0:19] sb_1__1__4_chanx_right_out;
  wire [0:19] sb_1__1__4_chany_bottom_out;
  wire [0:19] sb_1__1__4_chany_top_out;
  wire [0:0] sb_1__1__50_ccff_tail;
  wire [0:19] sb_1__1__50_chanx_left_out;
  wire [0:19] sb_1__1__50_chanx_right_out;
  wire [0:19] sb_1__1__50_chany_bottom_out;
  wire [0:19] sb_1__1__50_chany_top_out;
  wire [0:0] sb_1__1__51_ccff_tail;
  wire [0:19] sb_1__1__51_chanx_left_out;
  wire [0:19] sb_1__1__51_chanx_right_out;
  wire [0:19] sb_1__1__51_chany_bottom_out;
  wire [0:19] sb_1__1__51_chany_top_out;
  wire [0:0] sb_1__1__52_ccff_tail;
  wire [0:19] sb_1__1__52_chanx_left_out;
  wire [0:19] sb_1__1__52_chanx_right_out;
  wire [0:19] sb_1__1__52_chany_bottom_out;
  wire [0:19] sb_1__1__52_chany_top_out;
  wire [0:0] sb_1__1__53_ccff_tail;
  wire [0:19] sb_1__1__53_chanx_left_out;
  wire [0:19] sb_1__1__53_chanx_right_out;
  wire [0:19] sb_1__1__53_chany_bottom_out;
  wire [0:19] sb_1__1__53_chany_top_out;
  wire [0:0] sb_1__1__54_ccff_tail;
  wire [0:19] sb_1__1__54_chanx_left_out;
  wire [0:19] sb_1__1__54_chanx_right_out;
  wire [0:19] sb_1__1__54_chany_bottom_out;
  wire [0:19] sb_1__1__54_chany_top_out;
  wire [0:0] sb_1__1__55_ccff_tail;
  wire [0:19] sb_1__1__55_chanx_left_out;
  wire [0:19] sb_1__1__55_chanx_right_out;
  wire [0:19] sb_1__1__55_chany_bottom_out;
  wire [0:19] sb_1__1__55_chany_top_out;
  wire [0:0] sb_1__1__56_ccff_tail;
  wire [0:19] sb_1__1__56_chanx_left_out;
  wire [0:19] sb_1__1__56_chanx_right_out;
  wire [0:19] sb_1__1__56_chany_bottom_out;
  wire [0:19] sb_1__1__56_chany_top_out;
  wire [0:0] sb_1__1__57_ccff_tail;
  wire [0:19] sb_1__1__57_chanx_left_out;
  wire [0:19] sb_1__1__57_chanx_right_out;
  wire [0:19] sb_1__1__57_chany_bottom_out;
  wire [0:19] sb_1__1__57_chany_top_out;
  wire [0:0] sb_1__1__58_ccff_tail;
  wire [0:19] sb_1__1__58_chanx_left_out;
  wire [0:19] sb_1__1__58_chanx_right_out;
  wire [0:19] sb_1__1__58_chany_bottom_out;
  wire [0:19] sb_1__1__58_chany_top_out;
  wire [0:0] sb_1__1__59_ccff_tail;
  wire [0:19] sb_1__1__59_chanx_left_out;
  wire [0:19] sb_1__1__59_chanx_right_out;
  wire [0:19] sb_1__1__59_chany_bottom_out;
  wire [0:19] sb_1__1__59_chany_top_out;
  wire [0:0] sb_1__1__5_ccff_tail;
  wire [0:19] sb_1__1__5_chanx_left_out;
  wire [0:19] sb_1__1__5_chanx_right_out;
  wire [0:19] sb_1__1__5_chany_bottom_out;
  wire [0:19] sb_1__1__5_chany_top_out;
  wire [0:0] sb_1__1__60_ccff_tail;
  wire [0:19] sb_1__1__60_chanx_left_out;
  wire [0:19] sb_1__1__60_chanx_right_out;
  wire [0:19] sb_1__1__60_chany_bottom_out;
  wire [0:19] sb_1__1__60_chany_top_out;
  wire [0:0] sb_1__1__61_ccff_tail;
  wire [0:19] sb_1__1__61_chanx_left_out;
  wire [0:19] sb_1__1__61_chanx_right_out;
  wire [0:19] sb_1__1__61_chany_bottom_out;
  wire [0:19] sb_1__1__61_chany_top_out;
  wire [0:0] sb_1__1__62_ccff_tail;
  wire [0:19] sb_1__1__62_chanx_left_out;
  wire [0:19] sb_1__1__62_chanx_right_out;
  wire [0:19] sb_1__1__62_chany_bottom_out;
  wire [0:19] sb_1__1__62_chany_top_out;
  wire [0:0] sb_1__1__63_ccff_tail;
  wire [0:19] sb_1__1__63_chanx_left_out;
  wire [0:19] sb_1__1__63_chanx_right_out;
  wire [0:19] sb_1__1__63_chany_bottom_out;
  wire [0:19] sb_1__1__63_chany_top_out;
  wire [0:0] sb_1__1__64_ccff_tail;
  wire [0:19] sb_1__1__64_chanx_left_out;
  wire [0:19] sb_1__1__64_chanx_right_out;
  wire [0:19] sb_1__1__64_chany_bottom_out;
  wire [0:19] sb_1__1__64_chany_top_out;
  wire [0:0] sb_1__1__65_ccff_tail;
  wire [0:19] sb_1__1__65_chanx_left_out;
  wire [0:19] sb_1__1__65_chanx_right_out;
  wire [0:19] sb_1__1__65_chany_bottom_out;
  wire [0:19] sb_1__1__65_chany_top_out;
  wire [0:0] sb_1__1__66_ccff_tail;
  wire [0:19] sb_1__1__66_chanx_left_out;
  wire [0:19] sb_1__1__66_chanx_right_out;
  wire [0:19] sb_1__1__66_chany_bottom_out;
  wire [0:19] sb_1__1__66_chany_top_out;
  wire [0:0] sb_1__1__67_ccff_tail;
  wire [0:19] sb_1__1__67_chanx_left_out;
  wire [0:19] sb_1__1__67_chanx_right_out;
  wire [0:19] sb_1__1__67_chany_bottom_out;
  wire [0:19] sb_1__1__67_chany_top_out;
  wire [0:0] sb_1__1__68_ccff_tail;
  wire [0:19] sb_1__1__68_chanx_left_out;
  wire [0:19] sb_1__1__68_chanx_right_out;
  wire [0:19] sb_1__1__68_chany_bottom_out;
  wire [0:19] sb_1__1__68_chany_top_out;
  wire [0:0] sb_1__1__69_ccff_tail;
  wire [0:19] sb_1__1__69_chanx_left_out;
  wire [0:19] sb_1__1__69_chanx_right_out;
  wire [0:19] sb_1__1__69_chany_bottom_out;
  wire [0:19] sb_1__1__69_chany_top_out;
  wire [0:0] sb_1__1__6_ccff_tail;
  wire [0:19] sb_1__1__6_chanx_left_out;
  wire [0:19] sb_1__1__6_chanx_right_out;
  wire [0:19] sb_1__1__6_chany_bottom_out;
  wire [0:19] sb_1__1__6_chany_top_out;
  wire [0:0] sb_1__1__70_ccff_tail;
  wire [0:19] sb_1__1__70_chanx_left_out;
  wire [0:19] sb_1__1__70_chanx_right_out;
  wire [0:19] sb_1__1__70_chany_bottom_out;
  wire [0:19] sb_1__1__70_chany_top_out;
  wire [0:0] sb_1__1__71_ccff_tail;
  wire [0:19] sb_1__1__71_chanx_left_out;
  wire [0:19] sb_1__1__71_chanx_right_out;
  wire [0:19] sb_1__1__71_chany_bottom_out;
  wire [0:19] sb_1__1__71_chany_top_out;
  wire [0:0] sb_1__1__72_ccff_tail;
  wire [0:19] sb_1__1__72_chanx_left_out;
  wire [0:19] sb_1__1__72_chanx_right_out;
  wire [0:19] sb_1__1__72_chany_bottom_out;
  wire [0:19] sb_1__1__72_chany_top_out;
  wire [0:0] sb_1__1__73_ccff_tail;
  wire [0:19] sb_1__1__73_chanx_left_out;
  wire [0:19] sb_1__1__73_chanx_right_out;
  wire [0:19] sb_1__1__73_chany_bottom_out;
  wire [0:19] sb_1__1__73_chany_top_out;
  wire [0:0] sb_1__1__74_ccff_tail;
  wire [0:19] sb_1__1__74_chanx_left_out;
  wire [0:19] sb_1__1__74_chanx_right_out;
  wire [0:19] sb_1__1__74_chany_bottom_out;
  wire [0:19] sb_1__1__74_chany_top_out;
  wire [0:0] sb_1__1__75_ccff_tail;
  wire [0:19] sb_1__1__75_chanx_left_out;
  wire [0:19] sb_1__1__75_chanx_right_out;
  wire [0:19] sb_1__1__75_chany_bottom_out;
  wire [0:19] sb_1__1__75_chany_top_out;
  wire [0:0] sb_1__1__76_ccff_tail;
  wire [0:19] sb_1__1__76_chanx_left_out;
  wire [0:19] sb_1__1__76_chanx_right_out;
  wire [0:19] sb_1__1__76_chany_bottom_out;
  wire [0:19] sb_1__1__76_chany_top_out;
  wire [0:0] sb_1__1__7_ccff_tail;
  wire [0:19] sb_1__1__7_chanx_left_out;
  wire [0:19] sb_1__1__7_chanx_right_out;
  wire [0:19] sb_1__1__7_chany_bottom_out;
  wire [0:19] sb_1__1__7_chany_top_out;
  wire [0:0] sb_1__1__8_ccff_tail;
  wire [0:19] sb_1__1__8_chanx_left_out;
  wire [0:19] sb_1__1__8_chanx_right_out;
  wire [0:19] sb_1__1__8_chany_bottom_out;
  wire [0:19] sb_1__1__8_chany_top_out;
  wire [0:0] sb_1__1__9_ccff_tail;
  wire [0:19] sb_1__1__9_chanx_left_out;
  wire [0:19] sb_1__1__9_chanx_right_out;
  wire [0:19] sb_1__1__9_chany_bottom_out;
  wire [0:19] sb_1__1__9_chany_top_out;
  wire [0:0] sb_1__2__0_ccff_tail;
  wire [0:19] sb_1__2__0_chanx_left_out;
  wire [0:19] sb_1__2__0_chanx_right_out;
  wire [0:19] sb_1__2__0_chany_bottom_out;
  wire [0:19] sb_1__2__0_chany_top_out;
  wire [0:0] sb_1__2__10_ccff_tail;
  wire [0:19] sb_1__2__10_chanx_left_out;
  wire [0:19] sb_1__2__10_chanx_right_out;
  wire [0:19] sb_1__2__10_chany_bottom_out;
  wire [0:19] sb_1__2__10_chany_top_out;
  wire [0:0] sb_1__2__11_ccff_tail;
  wire [0:19] sb_1__2__11_chanx_left_out;
  wire [0:19] sb_1__2__11_chanx_right_out;
  wire [0:19] sb_1__2__11_chany_bottom_out;
  wire [0:19] sb_1__2__11_chany_top_out;
  wire [0:0] sb_1__2__1_ccff_tail;
  wire [0:19] sb_1__2__1_chanx_left_out;
  wire [0:19] sb_1__2__1_chanx_right_out;
  wire [0:19] sb_1__2__1_chany_bottom_out;
  wire [0:19] sb_1__2__1_chany_top_out;
  wire [0:0] sb_1__2__2_ccff_tail;
  wire [0:19] sb_1__2__2_chanx_left_out;
  wire [0:19] sb_1__2__2_chanx_right_out;
  wire [0:19] sb_1__2__2_chany_bottom_out;
  wire [0:19] sb_1__2__2_chany_top_out;
  wire [0:0] sb_1__2__3_ccff_tail;
  wire [0:19] sb_1__2__3_chanx_left_out;
  wire [0:19] sb_1__2__3_chanx_right_out;
  wire [0:19] sb_1__2__3_chany_bottom_out;
  wire [0:19] sb_1__2__3_chany_top_out;
  wire [0:0] sb_1__2__4_ccff_tail;
  wire [0:19] sb_1__2__4_chanx_left_out;
  wire [0:19] sb_1__2__4_chanx_right_out;
  wire [0:19] sb_1__2__4_chany_bottom_out;
  wire [0:19] sb_1__2__4_chany_top_out;
  wire [0:0] sb_1__2__5_ccff_tail;
  wire [0:19] sb_1__2__5_chanx_left_out;
  wire [0:19] sb_1__2__5_chanx_right_out;
  wire [0:19] sb_1__2__5_chany_bottom_out;
  wire [0:19] sb_1__2__5_chany_top_out;
  wire [0:0] sb_1__2__6_ccff_tail;
  wire [0:19] sb_1__2__6_chanx_left_out;
  wire [0:19] sb_1__2__6_chanx_right_out;
  wire [0:19] sb_1__2__6_chany_bottom_out;
  wire [0:19] sb_1__2__6_chany_top_out;
  wire [0:0] sb_1__2__7_ccff_tail;
  wire [0:19] sb_1__2__7_chanx_left_out;
  wire [0:19] sb_1__2__7_chanx_right_out;
  wire [0:19] sb_1__2__7_chany_bottom_out;
  wire [0:19] sb_1__2__7_chany_top_out;
  wire [0:0] sb_1__2__8_ccff_tail;
  wire [0:19] sb_1__2__8_chanx_left_out;
  wire [0:19] sb_1__2__8_chanx_right_out;
  wire [0:19] sb_1__2__8_chany_bottom_out;
  wire [0:19] sb_1__2__8_chany_top_out;
  wire [0:0] sb_1__2__9_ccff_tail;
  wire [0:19] sb_1__2__9_chanx_left_out;
  wire [0:19] sb_1__2__9_chanx_right_out;
  wire [0:19] sb_1__2__9_chany_bottom_out;
  wire [0:19] sb_1__2__9_chany_top_out;
  wire [0:0] sb_1__3__0_ccff_tail;
  wire [0:19] sb_1__3__0_chanx_left_out;
  wire [0:19] sb_1__3__0_chanx_right_out;
  wire [0:19] sb_1__3__0_chany_bottom_out;
  wire [0:19] sb_1__3__0_chany_top_out;
  wire [0:0] sb_1__3__10_ccff_tail;
  wire [0:19] sb_1__3__10_chanx_left_out;
  wire [0:19] sb_1__3__10_chanx_right_out;
  wire [0:19] sb_1__3__10_chany_bottom_out;
  wire [0:19] sb_1__3__10_chany_top_out;
  wire [0:0] sb_1__3__11_ccff_tail;
  wire [0:19] sb_1__3__11_chanx_left_out;
  wire [0:19] sb_1__3__11_chanx_right_out;
  wire [0:19] sb_1__3__11_chany_bottom_out;
  wire [0:19] sb_1__3__11_chany_top_out;
  wire [0:0] sb_1__3__1_ccff_tail;
  wire [0:19] sb_1__3__1_chanx_left_out;
  wire [0:19] sb_1__3__1_chanx_right_out;
  wire [0:19] sb_1__3__1_chany_bottom_out;
  wire [0:19] sb_1__3__1_chany_top_out;
  wire [0:0] sb_1__3__2_ccff_tail;
  wire [0:19] sb_1__3__2_chanx_left_out;
  wire [0:19] sb_1__3__2_chanx_right_out;
  wire [0:19] sb_1__3__2_chany_bottom_out;
  wire [0:19] sb_1__3__2_chany_top_out;
  wire [0:0] sb_1__3__3_ccff_tail;
  wire [0:19] sb_1__3__3_chanx_left_out;
  wire [0:19] sb_1__3__3_chanx_right_out;
  wire [0:19] sb_1__3__3_chany_bottom_out;
  wire [0:19] sb_1__3__3_chany_top_out;
  wire [0:0] sb_1__3__4_ccff_tail;
  wire [0:19] sb_1__3__4_chanx_left_out;
  wire [0:19] sb_1__3__4_chanx_right_out;
  wire [0:19] sb_1__3__4_chany_bottom_out;
  wire [0:19] sb_1__3__4_chany_top_out;
  wire [0:0] sb_1__3__5_ccff_tail;
  wire [0:19] sb_1__3__5_chanx_left_out;
  wire [0:19] sb_1__3__5_chanx_right_out;
  wire [0:19] sb_1__3__5_chany_bottom_out;
  wire [0:19] sb_1__3__5_chany_top_out;
  wire [0:0] sb_1__3__6_ccff_tail;
  wire [0:19] sb_1__3__6_chanx_left_out;
  wire [0:19] sb_1__3__6_chanx_right_out;
  wire [0:19] sb_1__3__6_chany_bottom_out;
  wire [0:19] sb_1__3__6_chany_top_out;
  wire [0:0] sb_1__3__7_ccff_tail;
  wire [0:19] sb_1__3__7_chanx_left_out;
  wire [0:19] sb_1__3__7_chanx_right_out;
  wire [0:19] sb_1__3__7_chany_bottom_out;
  wire [0:19] sb_1__3__7_chany_top_out;
  wire [0:0] sb_1__3__8_ccff_tail;
  wire [0:19] sb_1__3__8_chanx_left_out;
  wire [0:19] sb_1__3__8_chanx_right_out;
  wire [0:19] sb_1__3__8_chany_bottom_out;
  wire [0:19] sb_1__3__8_chany_top_out;
  wire [0:0] sb_1__3__9_ccff_tail;
  wire [0:19] sb_1__3__9_chanx_left_out;
  wire [0:19] sb_1__3__9_chanx_right_out;
  wire [0:19] sb_1__3__9_chany_bottom_out;
  wire [0:19] sb_1__3__9_chany_top_out;
  wire [0:0] sb_2__2__0_ccff_tail;
  wire [0:19] sb_2__2__0_chanx_left_out;
  wire [0:19] sb_2__2__0_chanx_right_out;
  wire [0:19] sb_2__2__0_chany_bottom_out;
  wire [0:19] sb_2__2__0_chany_top_out;
  wire [0:0] sb_2__2__1_ccff_tail;
  wire [0:19] sb_2__2__1_chanx_left_out;
  wire [0:19] sb_2__2__1_chanx_right_out;
  wire [0:19] sb_2__2__1_chany_bottom_out;
  wire [0:19] sb_2__2__1_chany_top_out;
  wire [0:0] sb_2__2__2_ccff_tail;
  wire [0:19] sb_2__2__2_chanx_left_out;
  wire [0:19] sb_2__2__2_chanx_right_out;
  wire [0:19] sb_2__2__2_chany_bottom_out;
  wire [0:19] sb_2__2__2_chany_top_out;
  wire [0:0] sb_2__2__3_ccff_tail;
  wire [0:19] sb_2__2__3_chanx_left_out;
  wire [0:19] sb_2__2__3_chanx_right_out;
  wire [0:19] sb_2__2__3_chany_bottom_out;
  wire [0:19] sb_2__2__3_chany_top_out;
  wire [0:0] sb_2__2__4_ccff_tail;
  wire [0:19] sb_2__2__4_chanx_left_out;
  wire [0:19] sb_2__2__4_chanx_right_out;
  wire [0:19] sb_2__2__4_chany_bottom_out;
  wire [0:19] sb_2__2__4_chany_top_out;
  wire [0:0] sb_2__2__5_ccff_tail;
  wire [0:19] sb_2__2__5_chanx_left_out;
  wire [0:19] sb_2__2__5_chanx_right_out;
  wire [0:19] sb_2__2__5_chany_bottom_out;
  wire [0:19] sb_2__2__5_chany_top_out;
  wire [0:0] sb_2__2__6_ccff_tail;
  wire [0:19] sb_2__2__6_chanx_left_out;
  wire [0:19] sb_2__2__6_chanx_right_out;
  wire [0:19] sb_2__2__6_chany_bottom_out;
  wire [0:19] sb_2__2__6_chany_top_out;
  wire [0:0] sb_2__2__7_ccff_tail;
  wire [0:19] sb_2__2__7_chanx_left_out;
  wire [0:19] sb_2__2__7_chanx_right_out;
  wire [0:19] sb_2__2__7_chany_bottom_out;
  wire [0:19] sb_2__2__7_chany_top_out;
  wire [0:0] sb_2__2__8_ccff_tail;
  wire [0:19] sb_2__2__8_chanx_left_out;
  wire [0:19] sb_2__2__8_chanx_right_out;
  wire [0:19] sb_2__2__8_chany_bottom_out;
  wire [0:19] sb_2__2__8_chany_top_out;
  wire [0:0] sb_2__2__9_ccff_tail;
  wire [0:19] sb_2__2__9_chanx_left_out;
  wire [0:19] sb_2__2__9_chanx_right_out;
  wire [0:19] sb_2__2__9_chany_bottom_out;
  wire [0:19] sb_2__2__9_chany_top_out;
  wire [0:0] sb_2__3__0_ccff_tail;
  wire [0:19] sb_2__3__0_chanx_left_out;
  wire [0:19] sb_2__3__0_chanx_right_out;
  wire [0:19] sb_2__3__0_chany_bottom_out;
  wire [0:19] sb_2__3__0_chany_top_out;
  wire [0:0] sb_2__3__1_ccff_tail;
  wire [0:19] sb_2__3__1_chanx_left_out;
  wire [0:19] sb_2__3__1_chanx_right_out;
  wire [0:19] sb_2__3__1_chany_bottom_out;
  wire [0:19] sb_2__3__1_chany_top_out;
  wire [0:0] sb_2__3__2_ccff_tail;
  wire [0:19] sb_2__3__2_chanx_left_out;
  wire [0:19] sb_2__3__2_chanx_right_out;
  wire [0:19] sb_2__3__2_chany_bottom_out;
  wire [0:19] sb_2__3__2_chany_top_out;
  wire [0:0] sb_2__3__3_ccff_tail;
  wire [0:19] sb_2__3__3_chanx_left_out;
  wire [0:19] sb_2__3__3_chanx_right_out;
  wire [0:19] sb_2__3__3_chany_bottom_out;
  wire [0:19] sb_2__3__3_chany_top_out;
  wire [0:0] sb_2__3__4_ccff_tail;
  wire [0:19] sb_2__3__4_chanx_left_out;
  wire [0:19] sb_2__3__4_chanx_right_out;
  wire [0:19] sb_2__3__4_chany_bottom_out;
  wire [0:19] sb_2__3__4_chany_top_out;
  wire [0:0] sb_2__3__5_ccff_tail;
  wire [0:19] sb_2__3__5_chanx_left_out;
  wire [0:19] sb_2__3__5_chanx_right_out;
  wire [0:19] sb_2__3__5_chany_bottom_out;
  wire [0:19] sb_2__3__5_chany_top_out;
  wire [0:0] sb_2__3__6_ccff_tail;
  wire [0:19] sb_2__3__6_chanx_left_out;
  wire [0:19] sb_2__3__6_chanx_right_out;
  wire [0:19] sb_2__3__6_chany_bottom_out;
  wire [0:19] sb_2__3__6_chany_top_out;
  wire [0:0] sb_2__3__7_ccff_tail;
  wire [0:19] sb_2__3__7_chanx_left_out;
  wire [0:19] sb_2__3__7_chanx_right_out;
  wire [0:19] sb_2__3__7_chany_bottom_out;
  wire [0:19] sb_2__3__7_chany_top_out;
  wire [0:0] sb_2__3__8_ccff_tail;
  wire [0:19] sb_2__3__8_chanx_left_out;
  wire [0:19] sb_2__3__8_chanx_right_out;
  wire [0:19] sb_2__3__8_chany_bottom_out;
  wire [0:19] sb_2__3__8_chany_top_out;
  wire [0:0] sb_2__3__9_ccff_tail;
  wire [0:19] sb_2__3__9_chanx_left_out;
  wire [0:19] sb_2__3__9_chanx_right_out;
  wire [0:19] sb_2__3__9_chany_bottom_out;
  wire [0:19] sb_2__3__9_chany_top_out;

  grid_clb
  grid_clb_1__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_84_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_0_ccff_tail)
  );


  grid_clb
  grid_clb_1__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_1_ccff_tail)
  );


  grid_clb
  grid_clb_1__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_85_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_2_ccff_tail)
  );


  grid_clb
  grid_clb_1__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_86_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_3_ccff_tail)
  );


  grid_clb
  grid_clb_1__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_87_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_4_ccff_tail)
  );


  grid_clb
  grid_clb_1__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_88_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_5_ccff_tail)
  );


  grid_clb
  grid_clb_1__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_89_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_6_ccff_tail)
  );


  grid_clb
  grid_clb_1__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_7_ccff_tail)
  );


  grid_clb
  grid_clb_1__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_90_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_8_ccff_tail)
  );


  grid_clb
  grid_clb_1__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_9_ccff_tail)
  );


  grid_clb
  grid_clb_2__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_91_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__10_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_10_ccff_tail)
  );


  grid_clb
  grid_clb_2__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__11_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_11_ccff_tail)
  );


  grid_clb
  grid_clb_2__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_92_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__12_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_12_ccff_tail)
  );


  grid_clb
  grid_clb_2__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_93_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__13_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_13_ccff_tail)
  );


  grid_clb
  grid_clb_2__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_94_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__14_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_14_ccff_tail)
  );


  grid_clb
  grid_clb_2__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_95_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__15_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_15_ccff_tail)
  );


  grid_clb
  grid_clb_2__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_96_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__16_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_16_ccff_tail)
  );


  grid_clb
  grid_clb_2__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__17_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_17_ccff_tail)
  );


  grid_clb
  grid_clb_2__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_97_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__18_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_18_ccff_tail)
  );


  grid_clb
  grid_clb_2__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_168_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__19_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_19_ccff_tail)
  );


  grid_clb
  grid_clb_3__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_98_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__20_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_20_ccff_tail)
  );


  grid_clb
  grid_clb_3__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__21_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_21_ccff_tail)
  );


  grid_clb
  grid_clb_3__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_99_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__22_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_22_ccff_tail)
  );


  grid_clb
  grid_clb_3__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_100_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__23_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_23_ccff_tail)
  );


  grid_clb
  grid_clb_3__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_101_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__24_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_24_ccff_tail)
  );


  grid_clb
  grid_clb_3__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_102_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__25_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_25_ccff_tail)
  );


  grid_clb
  grid_clb_3__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_103_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__26_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_26_ccff_tail)
  );


  grid_clb
  grid_clb_3__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__27_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_27_ccff_tail)
  );


  grid_clb
  grid_clb_3__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_104_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__28_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_28_ccff_tail)
  );


  grid_clb
  grid_clb_3__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_169_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__29_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_29_ccff_tail)
  );


  grid_clb
  grid_clb_4__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_105_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__30_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_30_ccff_tail)
  );


  grid_clb
  grid_clb_4__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__31_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_31_ccff_tail)
  );


  grid_clb
  grid_clb_4__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_106_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__32_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_32_ccff_tail)
  );


  grid_clb
  grid_clb_4__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_107_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__33_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_33_ccff_tail)
  );


  grid_clb
  grid_clb_4__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_108_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__34_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_34_ccff_tail)
  );


  grid_clb
  grid_clb_4__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_109_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__35_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_35_ccff_tail)
  );


  grid_clb
  grid_clb_4__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_110_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__36_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_36_ccff_tail)
  );


  grid_clb
  grid_clb_4__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__37_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_37_ccff_tail)
  );


  grid_clb
  grid_clb_4__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_111_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__38_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_38_ccff_tail)
  );


  grid_clb
  grid_clb_4__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_170_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__39_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_39_ccff_tail)
  );


  grid_clb
  grid_clb_5__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_112_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_28_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__40_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_40_ccff_tail)
  );


  grid_clb
  grid_clb_5__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__41_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_41_ccff_tail)
  );


  grid_clb
  grid_clb_5__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_113_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_29_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__42_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_42_ccff_tail)
  );


  grid_clb
  grid_clb_5__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_114_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_30_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__43_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_43_ccff_tail)
  );


  grid_clb
  grid_clb_5__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_115_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_31_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__44_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_44_ccff_tail)
  );


  grid_clb
  grid_clb_5__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_116_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_32_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__45_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_45_ccff_tail)
  );


  grid_clb
  grid_clb_5__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_117_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_33_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__46_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_46_ccff_tail)
  );


  grid_clb
  grid_clb_5__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__47_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_47_ccff_tail)
  );


  grid_clb
  grid_clb_5__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_118_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_34_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__48_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_48_ccff_tail)
  );


  grid_clb
  grid_clb_5__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_171_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__49_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_49_ccff_tail)
  );


  grid_clb
  grid_clb_6__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_119_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_35_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__50_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_50_ccff_tail)
  );


  grid_clb
  grid_clb_6__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__51_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_51_ccff_tail)
  );


  grid_clb
  grid_clb_6__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_120_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_36_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__52_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_52_ccff_tail)
  );


  grid_clb
  grid_clb_6__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_121_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_37_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__53_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_53_ccff_tail)
  );


  grid_clb
  grid_clb_6__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_122_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_38_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__54_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_54_ccff_tail)
  );


  grid_clb
  grid_clb_6__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_123_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_39_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__55_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_55_ccff_tail)
  );


  grid_clb
  grid_clb_6__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_124_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_40_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__56_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_56_ccff_tail)
  );


  grid_clb
  grid_clb_6__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__57_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_57_ccff_tail)
  );


  grid_clb
  grid_clb_6__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_125_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_41_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__58_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_58_ccff_tail)
  );


  grid_clb
  grid_clb_6__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_172_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__59_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_59_ccff_tail)
  );


  grid_clb
  grid_clb_7__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_126_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_42_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__60_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_60_ccff_tail)
  );


  grid_clb
  grid_clb_7__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__61_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_61_ccff_tail)
  );


  grid_clb
  grid_clb_7__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_127_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_43_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__62_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_62_ccff_tail)
  );


  grid_clb
  grid_clb_7__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_128_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_44_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__63_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_63_ccff_tail)
  );


  grid_clb
  grid_clb_7__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_129_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_45_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__64_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_64_ccff_tail)
  );


  grid_clb
  grid_clb_7__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_130_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_46_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__65_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_65_ccff_tail)
  );


  grid_clb
  grid_clb_7__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_131_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_47_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__66_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_66_ccff_tail)
  );


  grid_clb
  grid_clb_7__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__67_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_67_ccff_tail)
  );


  grid_clb
  grid_clb_7__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_132_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_48_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__68_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_68_ccff_tail)
  );


  grid_clb
  grid_clb_7__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_173_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__69_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_69_ccff_tail)
  );


  grid_clb
  grid_clb_8__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_133_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_49_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__70_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_70_ccff_tail)
  );


  grid_clb
  grid_clb_8__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__71_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_71_ccff_tail)
  );


  grid_clb
  grid_clb_8__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_134_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_50_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__72_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_72_ccff_tail)
  );


  grid_clb
  grid_clb_8__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_135_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_51_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__73_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_73_ccff_tail)
  );


  grid_clb
  grid_clb_8__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_136_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_52_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__74_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_74_ccff_tail)
  );


  grid_clb
  grid_clb_8__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_137_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_53_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__75_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_75_ccff_tail)
  );


  grid_clb
  grid_clb_8__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_138_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_54_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__76_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_76_ccff_tail)
  );


  grid_clb
  grid_clb_8__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__77_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_77_ccff_tail)
  );


  grid_clb
  grid_clb_8__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_139_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_55_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__78_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_78_ccff_tail)
  );


  grid_clb
  grid_clb_8__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_174_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__79_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_79_ccff_tail)
  );


  grid_clb
  grid_clb_9__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_140_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_56_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__80_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_80_ccff_tail)
  );


  grid_clb
  grid_clb_9__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__81_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_81_ccff_tail)
  );


  grid_clb
  grid_clb_9__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_141_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_57_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__82_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_82_ccff_tail)
  );


  grid_clb
  grid_clb_9__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_142_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_58_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__83_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_83_ccff_tail)
  );


  grid_clb
  grid_clb_9__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_143_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_59_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__84_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_84_ccff_tail)
  );


  grid_clb
  grid_clb_9__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_144_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_60_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__85_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_85_ccff_tail)
  );


  grid_clb
  grid_clb_9__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_145_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_61_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__86_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_86_ccff_tail)
  );


  grid_clb
  grid_clb_9__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__87_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_87_ccff_tail)
  );


  grid_clb
  grid_clb_9__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_146_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_62_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__88_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_88_ccff_tail)
  );


  grid_clb
  grid_clb_9__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_175_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__89_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_89_ccff_tail)
  );


  grid_clb
  grid_clb_10__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_147_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_63_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__90_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_90_ccff_tail)
  );


  grid_clb
  grid_clb_10__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__91_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_91_ccff_tail)
  );


  grid_clb
  grid_clb_10__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_148_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_64_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__92_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_92_ccff_tail)
  );


  grid_clb
  grid_clb_10__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_149_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_65_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__93_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_93_ccff_tail)
  );


  grid_clb
  grid_clb_10__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_150_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_66_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__94_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_94_ccff_tail)
  );


  grid_clb
  grid_clb_10__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_151_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_67_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__95_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_95_ccff_tail)
  );


  grid_clb
  grid_clb_10__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_152_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_68_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__96_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_96_ccff_tail)
  );


  grid_clb
  grid_clb_10__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__97_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_97_ccff_tail)
  );


  grid_clb
  grid_clb_10__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_153_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_69_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__98_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_98_ccff_tail)
  );


  grid_clb
  grid_clb_10__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_176_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_10__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__99_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_99_ccff_tail)
  );


  grid_clb
  grid_clb_11__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_154_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_70_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__100_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_100_ccff_tail)
  );


  grid_clb
  grid_clb_11__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__101_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_101_ccff_tail)
  );


  grid_clb
  grid_clb_11__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_155_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_71_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__102_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_102_ccff_tail)
  );


  grid_clb
  grid_clb_11__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_156_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_72_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__103_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_103_ccff_tail)
  );


  grid_clb
  grid_clb_11__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_157_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_73_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__104_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_104_ccff_tail)
  );


  grid_clb
  grid_clb_11__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_158_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_74_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__105_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_105_ccff_tail)
  );


  grid_clb
  grid_clb_11__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_159_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_75_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__106_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_106_ccff_tail)
  );


  grid_clb
  grid_clb_11__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__107_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_107_ccff_tail)
  );


  grid_clb
  grid_clb_11__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_160_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_76_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__108_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_108_ccff_tail)
  );


  grid_clb
  grid_clb_11__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_177_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_11__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(cby_1__1__109_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_109_ccff_tail)
  );


  grid_clb
  grid_clb_12__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_161_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_77_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_11_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_110_ccff_tail)
  );


  grid_clb
  grid_clb_12__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_10_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_111_ccff_tail)
  );


  grid_clb
  grid_clb_12__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_162_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_78_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_112_ccff_tail)
  );


  grid_clb
  grid_clb_12__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_163_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_79_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_113_ccff_tail)
  );


  grid_clb
  grid_clb_12__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_164_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_80_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_114_ccff_tail)
  );


  grid_clb
  grid_clb_12__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_165_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_81_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_115_ccff_tail)
  );


  grid_clb
  grid_clb_12__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_166_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_82_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_116_ccff_tail)
  );


  grid_clb
  grid_clb_12__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_117_ccff_tail)
  );


  grid_clb
  grid_clb_12__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_167_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_83_out),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_118_ccff_tail)
  );


  grid_clb
  grid_clb_12__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .Test_en(Test_en),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_178_out),
    .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_12__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .left_width_0_height_0_subtile_0__pin_reset_0_(reset),
    .left_width_0_height_0_subtile_0__pin_clk_0_(clk),
    .ccff_head(grid_io_right_right_0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .ccff_tail(grid_clb_119_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_1__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_0_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_1__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_1_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_3__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_2_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_3__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_3_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_5__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_4_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_5__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_5_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_7__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_6_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_7__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_7_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_9__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_8_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_9__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_9_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_11__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(grid_io_right_right_9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_10_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_11__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(grid_io_right_right_2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_11_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_1__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[0]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[0]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[0]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__0_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_0_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_2__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[1]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[1]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[1]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__1_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_1_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_3__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[2]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[2]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[2]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__2_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_2_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_4__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[3]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[3]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[3]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__3_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_3_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_5__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[4]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[4]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[4]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__4_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_4_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_6__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[5]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[5]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[5]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__5_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_5_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_7__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[6]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[6]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[6]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__6_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_6_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_8__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[7]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[7]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[7]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__7_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_7_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_9__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[8]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[8]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[8]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__8_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_8_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_10__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[9]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[9]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[9]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__9_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_9_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_11__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[10]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[10]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[10]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__10_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_10_ccff_tail)
  );


  grid_io_top_top
  grid_io_top_top_12__13_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[11]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[11]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[11]),
    .bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cbx_1__12__11_ccff_tail),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_11_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__12_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[12]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[12]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[12]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__9_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_0_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__11_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[13]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[13]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[13]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__8_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_1_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__10_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[14]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[14]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[14]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__3__1_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_2_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__9_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[15]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[15]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[15]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__7_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_3_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__8_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[16]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[16]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[16]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__6_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_4_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__7_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[17]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[17]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[17]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__5_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_5_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__6_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[18]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[18]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[18]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__4_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_6_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__5_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[19]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[19]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[19]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__3_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_7_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__4_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[20]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[20]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[20]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__2_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_8_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__3_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[21]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[21]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[21]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__3__0_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_9_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__2_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[22]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[22]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[22]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__1_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_10_ccff_tail)
  );


  grid_io_right_right
  grid_io_right_right_13__1_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[23]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[23]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[23]),
    .left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_12__1__0_ccff_tail),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_11_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_12__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[24:32]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[24:32]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[24:32]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__11_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_0_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_11__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[33:41]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[33:41]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[33:41]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__10_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_1_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_10__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[42:50]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[42:50]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[42:50]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_2_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_9__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[51:59]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[51:59]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[51:59]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_3_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_8__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[60:68]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[60:68]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[60:68]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_4_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_7__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[69:77]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[69:77]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[69:77]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_5_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_6__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[78:86]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[78:86]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[78:86]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_6_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_5__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[87:95]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[87:95]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[87:95]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_7_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_4__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[96:104]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[96:104]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[96:104]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_8_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_3__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[105:113]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[105:113]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[105:113]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_9_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_2__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[114:122]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[114:122]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[114:122]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_10_ccff_tail)
  );


  grid_io_bottom_bottom
  grid_io_bottom_bottom_1__0_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[123:131]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[123:131]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[123:131]),
    .top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_head(cbx_1__0__0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_11_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__1_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[132]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[132]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[132]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__0_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_0_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__2_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[133]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[133]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[133]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__1_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_1_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__3_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[134]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[134]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[134]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__2_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_2_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__4_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[135]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[135]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[135]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__3_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_3_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__5_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[136]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[136]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[136]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__4_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_4_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__6_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[137]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[137]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[137]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__5_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_5_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__7_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[138]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[138]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[138]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__6_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_6_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__8_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[139]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[139]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[139]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__7_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_7_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__9_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[140]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[140]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[140]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__8_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_8_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__10_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[141]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[141]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[141]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__9_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_9_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__11_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[142]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[142]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[142]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__10_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_10_ccff_tail)
  );


  grid_io_left_left
  grid_io_left_left_0__12_
  (
    .IO_ISOL_N(IO_ISOL_N),
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[143]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[143]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[143]),
    .right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_head(cby_0__1__11_ccff_tail),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_11_ccff_tail)
  );


  sb_0__0_
  sb_0__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_0_ccff_tail),
    .chany_top_out(sb_0__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
    .ccff_tail(sb_0__0__0_ccff_tail)
  );


  sb_0__1_
  sb_0__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_1_ccff_tail),
    .chany_top_out(sb_0__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__0_ccff_tail)
  );


  sb_0__1_
  sb_0__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_2_ccff_tail),
    .chany_top_out(sb_0__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__1_ccff_tail)
  );


  sb_0__1_
  sb_0__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_4_ccff_tail),
    .chany_top_out(sb_0__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__2_ccff_tail)
  );


  sb_0__1_
  sb_0__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_5_ccff_tail),
    .chany_top_out(sb_0__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__3_ccff_tail)
  );


  sb_0__1_
  sb_0__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_6_ccff_tail),
    .chany_top_out(sb_0__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__4_ccff_tail)
  );


  sb_0__1_
  sb_0__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_7_ccff_tail),
    .chany_top_out(sb_0__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__5_ccff_tail)
  );


  sb_0__1_
  sb_0__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_8_ccff_tail),
    .chany_top_out(sb_0__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__6_ccff_tail)
  );


  sb_0__1_
  sb_0__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_9_ccff_tail),
    .chany_top_out(sb_0__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__7_ccff_tail)
  );


  sb_0__1_
  sb_0__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__11_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__10_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_11_ccff_tail),
    .chany_top_out(sb_0__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__8_ccff_tail)
  );


  sb_0__3_
  sb_0__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__3__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_3_ccff_tail),
    .chany_top_out(sb_0__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__3__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__3__0_ccff_tail)
  );


  sb_0__3_
  sb_0__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_0__1__10_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__3__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_0__1__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_10_ccff_tail),
    .chany_top_out(sb_0__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__3__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__3__1_ccff_tail)
  );


  sb_0__12_
  sb_0__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__0_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__11_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_top_top_0_ccff_tail),
    .chanx_right_out(sb_0__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__12__0_ccff_tail)
  );


  sb_1__0_
  sb_1__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_11_ccff_tail),
    .chany_top_out(sb_1__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__0_ccff_tail)
  );


  sb_1__0_
  sb_2__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_10_ccff_tail),
    .chany_top_out(sb_1__0__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__1_ccff_tail)
  );


  sb_1__0_
  sb_3__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_9_ccff_tail),
    .chany_top_out(sb_1__0__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__2_ccff_tail)
  );


  sb_1__0_
  sb_4__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_8_ccff_tail),
    .chany_top_out(sb_1__0__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__3_ccff_tail)
  );


  sb_1__0_
  sb_5__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_7_ccff_tail),
    .chany_top_out(sb_1__0__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__4_ccff_tail)
  );


  sb_1__0_
  sb_6__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_6_ccff_tail),
    .chany_top_out(sb_1__0__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__5_ccff_tail)
  );


  sb_1__0_
  sb_7__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__60_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_5_ccff_tail),
    .chany_top_out(sb_1__0__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__6_ccff_tail)
  );


  sb_1__0_
  sb_8__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__70_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_4_ccff_tail),
    .chany_top_out(sb_1__0__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__7_ccff_tail)
  );


  sb_1__0_
  sb_9__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__80_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_3_ccff_tail),
    .chany_top_out(sb_1__0__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__8_ccff_tail)
  );


  sb_1__0_
  sb_10__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__90_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_2_ccff_tail),
    .chany_top_out(sb_1__0__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__9_ccff_tail)
  );


  sb_1__0_
  sb_11__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__100_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_1_ccff_tail),
    .chany_top_out(sb_1__0__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__10_ccff_tail)
  );


  sb_1__1_
  sb_1__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__0_ccff_tail),
    .chany_top_out(sb_1__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__0_ccff_tail)
  );


  sb_1__1_
  sb_1__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__2_ccff_tail),
    .chany_top_out(sb_1__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__1_ccff_tail)
  );


  sb_1__1_
  sb_1__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__3_ccff_tail),
    .chany_top_out(sb_1__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__2_ccff_tail)
  );


  sb_1__1_
  sb_1__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__4_ccff_tail),
    .chany_top_out(sb_1__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__3_ccff_tail)
  );


  sb_1__1_
  sb_1__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__5_ccff_tail),
    .chany_top_out(sb_1__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__4_ccff_tail)
  );


  sb_1__1_
  sb_1__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__6_ccff_tail),
    .chany_top_out(sb_1__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__5_ccff_tail)
  );


  sb_1__1_
  sb_1__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__8_ccff_tail),
    .chany_top_out(sb_1__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__6_ccff_tail)
  );


  sb_1__1_
  sb_2__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__9_ccff_tail),
    .chany_top_out(sb_1__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__7_ccff_tail)
  );


  sb_1__1_
  sb_2__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__11_ccff_tail),
    .chany_top_out(sb_1__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__8_ccff_tail)
  );


  sb_1__1_
  sb_2__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__12_ccff_tail),
    .chany_top_out(sb_1__1__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__9_ccff_tail)
  );


  sb_1__1_
  sb_2__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__13_ccff_tail),
    .chany_top_out(sb_1__1__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__10_ccff_tail)
  );


  sb_1__1_
  sb_2__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__14_ccff_tail),
    .chany_top_out(sb_1__1__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__11_ccff_tail)
  );


  sb_1__1_
  sb_2__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__15_ccff_tail),
    .chany_top_out(sb_1__1__12_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__12_ccff_tail)
  );


  sb_1__1_
  sb_2__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__17_ccff_tail),
    .chany_top_out(sb_1__1__13_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__13_ccff_tail)
  );


  sb_1__1_
  sb_3__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__18_ccff_tail),
    .chany_top_out(sb_1__1__14_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__14_ccff_tail)
  );


  sb_1__1_
  sb_3__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__20_ccff_tail),
    .chany_top_out(sb_1__1__15_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__15_ccff_tail)
  );


  sb_1__1_
  sb_3__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__21_ccff_tail),
    .chany_top_out(sb_1__1__16_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__16_ccff_tail)
  );


  sb_1__1_
  sb_3__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__22_ccff_tail),
    .chany_top_out(sb_1__1__17_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__17_ccff_tail)
  );


  sb_1__1_
  sb_3__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__23_ccff_tail),
    .chany_top_out(sb_1__1__18_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__18_ccff_tail)
  );


  sb_1__1_
  sb_3__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__24_ccff_tail),
    .chany_top_out(sb_1__1__19_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__19_ccff_tail)
  );


  sb_1__1_
  sb_3__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__26_ccff_tail),
    .chany_top_out(sb_1__1__20_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__20_ccff_tail)
  );


  sb_1__1_
  sb_4__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__27_ccff_tail),
    .chany_top_out(sb_1__1__21_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__21_ccff_tail)
  );


  sb_1__1_
  sb_4__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__29_ccff_tail),
    .chany_top_out(sb_1__1__22_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__22_ccff_tail)
  );


  sb_1__1_
  sb_4__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__30_ccff_tail),
    .chany_top_out(sb_1__1__23_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__23_ccff_tail)
  );


  sb_1__1_
  sb_4__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__31_ccff_tail),
    .chany_top_out(sb_1__1__24_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__24_ccff_tail)
  );


  sb_1__1_
  sb_4__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__32_ccff_tail),
    .chany_top_out(sb_1__1__25_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__25_ccff_tail)
  );


  sb_1__1_
  sb_4__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__33_ccff_tail),
    .chany_top_out(sb_1__1__26_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__26_ccff_tail)
  );


  sb_1__1_
  sb_4__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__35_ccff_tail),
    .chany_top_out(sb_1__1__27_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__27_ccff_tail)
  );


  sb_1__1_
  sb_5__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__36_ccff_tail),
    .chany_top_out(sb_1__1__28_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__28_ccff_tail)
  );


  sb_1__1_
  sb_5__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__38_ccff_tail),
    .chany_top_out(sb_1__1__29_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__29_ccff_tail)
  );


  sb_1__1_
  sb_5__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__39_ccff_tail),
    .chany_top_out(sb_1__1__30_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__30_ccff_tail)
  );


  sb_1__1_
  sb_5__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__40_ccff_tail),
    .chany_top_out(sb_1__1__31_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__31_ccff_tail)
  );


  sb_1__1_
  sb_5__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__41_ccff_tail),
    .chany_top_out(sb_1__1__32_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__32_ccff_tail)
  );


  sb_1__1_
  sb_5__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__42_ccff_tail),
    .chany_top_out(sb_1__1__33_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__33_ccff_tail)
  );


  sb_1__1_
  sb_5__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__44_ccff_tail),
    .chany_top_out(sb_1__1__34_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__34_ccff_tail)
  );


  sb_1__1_
  sb_6__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__45_ccff_tail),
    .chany_top_out(sb_1__1__35_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__35_ccff_tail)
  );


  sb_1__1_
  sb_6__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__56_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__47_ccff_tail),
    .chany_top_out(sb_1__1__36_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__36_ccff_tail)
  );


  sb_1__1_
  sb_6__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__57_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__48_ccff_tail),
    .chany_top_out(sb_1__1__37_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__37_ccff_tail)
  );


  sb_1__1_
  sb_6__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__58_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__49_ccff_tail),
    .chany_top_out(sb_1__1__38_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__38_ccff_tail)
  );


  sb_1__1_
  sb_6__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__56_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__59_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__50_ccff_tail),
    .chany_top_out(sb_1__1__39_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__39_ccff_tail)
  );


  sb_1__1_
  sb_6__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__57_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__60_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__56_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__51_ccff_tail),
    .chany_top_out(sb_1__1__40_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__40_ccff_tail)
  );


  sb_1__1_
  sb_6__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__59_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__62_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__58_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__53_ccff_tail),
    .chany_top_out(sb_1__1__41_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__41_ccff_tail)
  );


  sb_1__1_
  sb_7__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__61_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__63_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__60_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__54_ccff_tail),
    .chany_top_out(sb_1__1__42_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__42_ccff_tail)
  );


  sb_1__1_
  sb_7__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__63_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__65_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__62_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__56_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__56_ccff_tail),
    .chany_top_out(sb_1__1__43_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__43_ccff_tail)
  );


  sb_1__1_
  sb_7__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__64_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__66_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__63_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__57_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__57_ccff_tail),
    .chany_top_out(sb_1__1__44_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__44_ccff_tail)
  );


  sb_1__1_
  sb_7__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__65_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__67_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__64_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__58_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__58_ccff_tail),
    .chany_top_out(sb_1__1__45_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__45_ccff_tail)
  );


  sb_1__1_
  sb_7__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__66_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__68_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__65_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__59_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__59_ccff_tail),
    .chany_top_out(sb_1__1__46_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__46_ccff_tail)
  );


  sb_1__1_
  sb_7__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__67_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__69_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__66_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__60_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__60_ccff_tail),
    .chany_top_out(sb_1__1__47_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__47_ccff_tail)
  );


  sb_1__1_
  sb_7__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__69_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__71_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__68_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__62_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__62_ccff_tail),
    .chany_top_out(sb_1__1__48_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__48_ccff_tail)
  );


  sb_1__1_
  sb_8__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__71_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__72_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__70_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__63_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__63_ccff_tail),
    .chany_top_out(sb_1__1__49_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__49_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__49_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__49_ccff_tail)
  );


  sb_1__1_
  sb_8__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__73_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__74_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__72_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__65_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__65_ccff_tail),
    .chany_top_out(sb_1__1__50_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__50_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__50_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__50_ccff_tail)
  );


  sb_1__1_
  sb_8__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__74_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__75_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__73_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__66_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__66_ccff_tail),
    .chany_top_out(sb_1__1__51_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__51_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__51_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__51_ccff_tail)
  );


  sb_1__1_
  sb_8__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__75_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__76_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__74_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__67_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__67_ccff_tail),
    .chany_top_out(sb_1__1__52_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__52_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__52_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__52_ccff_tail)
  );


  sb_1__1_
  sb_8__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__76_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__77_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__75_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__68_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__68_ccff_tail),
    .chany_top_out(sb_1__1__53_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__53_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__53_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__53_ccff_tail)
  );


  sb_1__1_
  sb_8__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__77_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__78_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__76_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__69_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__69_ccff_tail),
    .chany_top_out(sb_1__1__54_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__54_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__54_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__54_ccff_tail)
  );


  sb_1__1_
  sb_8__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__79_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__80_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__78_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__71_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__71_ccff_tail),
    .chany_top_out(sb_1__1__55_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__55_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__55_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__55_ccff_tail)
  );


  sb_1__1_
  sb_9__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__81_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__81_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__80_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__72_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__72_ccff_tail),
    .chany_top_out(sb_1__1__56_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__56_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__56_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__56_ccff_tail)
  );


  sb_1__1_
  sb_9__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__83_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__83_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__82_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__74_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__74_ccff_tail),
    .chany_top_out(sb_1__1__57_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__57_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__57_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__57_ccff_tail)
  );


  sb_1__1_
  sb_9__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__84_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__84_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__83_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__75_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__75_ccff_tail),
    .chany_top_out(sb_1__1__58_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__58_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__58_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__58_ccff_tail)
  );


  sb_1__1_
  sb_9__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__85_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__85_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__84_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__76_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__76_ccff_tail),
    .chany_top_out(sb_1__1__59_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__59_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__59_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__59_ccff_tail)
  );


  sb_1__1_
  sb_9__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__86_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__86_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__85_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__77_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__77_ccff_tail),
    .chany_top_out(sb_1__1__60_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__60_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__60_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__60_ccff_tail)
  );


  sb_1__1_
  sb_9__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__87_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__87_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__86_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__78_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__78_ccff_tail),
    .chany_top_out(sb_1__1__61_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__61_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__61_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__61_ccff_tail)
  );


  sb_1__1_
  sb_9__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__89_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__89_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__88_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__80_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__80_ccff_tail),
    .chany_top_out(sb_1__1__62_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__62_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__62_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__62_ccff_tail)
  );


  sb_1__1_
  sb_10__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__91_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__90_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__90_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__81_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__81_ccff_tail),
    .chany_top_out(sb_1__1__63_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__63_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__63_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__63_ccff_tail)
  );


  sb_1__1_
  sb_10__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__93_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__92_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__92_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__83_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__83_ccff_tail),
    .chany_top_out(sb_1__1__64_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__64_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__64_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__64_ccff_tail)
  );


  sb_1__1_
  sb_10__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__94_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__93_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__93_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__84_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__84_ccff_tail),
    .chany_top_out(sb_1__1__65_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__65_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__65_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__65_ccff_tail)
  );


  sb_1__1_
  sb_10__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__95_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__94_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__94_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__85_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__85_ccff_tail),
    .chany_top_out(sb_1__1__66_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__66_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__66_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__66_ccff_tail)
  );


  sb_1__1_
  sb_10__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__96_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__95_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__95_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__86_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__86_ccff_tail),
    .chany_top_out(sb_1__1__67_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__67_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__67_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__67_ccff_tail)
  );


  sb_1__1_
  sb_10__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__97_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__96_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__96_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__87_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__87_ccff_tail),
    .chany_top_out(sb_1__1__68_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__68_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__68_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__68_ccff_tail)
  );


  sb_1__1_
  sb_10__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__99_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__98_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__98_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__89_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__89_ccff_tail),
    .chany_top_out(sb_1__1__69_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__69_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__69_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__69_ccff_tail)
  );


  sb_1__1_
  sb_11__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__101_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__99_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__100_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__90_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__90_ccff_tail),
    .chany_top_out(sb_1__1__70_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__70_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__70_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__70_ccff_tail)
  );


  sb_1__1_
  sb_11__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__103_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__101_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__102_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__92_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__92_ccff_tail),
    .chany_top_out(sb_1__1__71_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__71_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__71_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__71_ccff_tail)
  );


  sb_1__1_
  sb_11__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__104_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__102_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__103_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__93_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__93_ccff_tail),
    .chany_top_out(sb_1__1__72_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__72_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__72_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__72_ccff_tail)
  );


  sb_1__1_
  sb_11__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__105_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__103_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__104_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__94_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__94_ccff_tail),
    .chany_top_out(sb_1__1__73_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__73_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__73_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__73_ccff_tail)
  );


  sb_1__1_
  sb_11__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__106_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__104_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__105_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__95_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__95_ccff_tail),
    .chany_top_out(sb_1__1__74_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__74_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__74_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__74_ccff_tail)
  );


  sb_1__1_
  sb_11__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__107_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__105_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__106_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__96_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__96_ccff_tail),
    .chany_top_out(sb_1__1__75_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__75_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__75_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__75_ccff_tail)
  );


  sb_1__1_
  sb_11__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__109_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__107_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__108_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__98_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__98_ccff_tail),
    .chany_top_out(sb_1__1__76_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__76_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__76_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__76_ccff_tail)
  );


  sb_1__2_
  sb_1__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__0_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__1_ccff_tail),
    .chany_top_out(sb_1__2__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__0_ccff_tail)
  );


  sb_1__2_
  sb_1__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__1_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__7_ccff_tail),
    .chany_top_out(sb_1__2__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__1_ccff_tail)
  );


  sb_1__2_
  sb_3__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__2_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__19_ccff_tail),
    .chany_top_out(sb_1__2__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__2_ccff_tail)
  );


  sb_1__2_
  sb_3__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__3_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__25_ccff_tail),
    .chany_top_out(sb_1__2__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__3_ccff_tail)
  );


  sb_1__2_
  sb_5__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__4_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__37_ccff_tail),
    .chany_top_out(sb_1__2__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__4_ccff_tail)
  );


  sb_1__2_
  sb_5__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__5_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__43_ccff_tail),
    .chany_top_out(sb_1__2__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__5_ccff_tail)
  );


  sb_1__2_
  sb_7__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__6_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__64_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__61_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__55_ccff_tail),
    .chany_top_out(sb_1__2__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__6_ccff_tail)
  );


  sb_1__2_
  sb_7__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__7_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__70_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__67_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__61_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__61_ccff_tail),
    .chany_top_out(sb_1__2__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__7_ccff_tail)
  );


  sb_1__2_
  sb_9__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__8_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__82_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__81_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__73_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__73_ccff_tail),
    .chany_top_out(sb_1__2__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__8_ccff_tail)
  );


  sb_1__2_
  sb_9__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__9_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__88_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__87_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__79_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__79_ccff_tail),
    .chany_top_out(sb_1__2__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__9_ccff_tail)
  );


  sb_1__2_
  sb_11__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__10_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__100_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__101_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__91_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__91_ccff_tail),
    .chany_top_out(sb_1__2__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__10_ccff_tail)
  );


  sb_1__2_
  sb_11__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__3__11_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__106_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__107_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__97_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__97_ccff_tail),
    .chany_top_out(sb_1__2__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__11_ccff_tail)
  );


  sb_1__3_
  sb_1__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__0_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__0_ccff_tail),
    .chany_top_out(sb_1__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__0_ccff_tail)
  );


  sb_1__3_
  sb_1__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__1_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__1_ccff_tail),
    .chany_top_out(sb_1__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__1_ccff_tail)
  );


  sb_1__3_
  sb_3__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__2_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__2_ccff_tail),
    .chany_top_out(sb_1__3__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__2_ccff_tail)
  );


  sb_1__3_
  sb_3__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__3_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__3_ccff_tail),
    .chany_top_out(sb_1__3__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__3_ccff_tail)
  );


  sb_1__3_
  sb_5__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__4_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__4_ccff_tail),
    .chany_top_out(sb_1__3__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__4_ccff_tail)
  );


  sb_1__3_
  sb_5__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__5_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__5_ccff_tail),
    .chany_top_out(sb_1__3__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__5_ccff_tail)
  );


  sb_1__3_
  sb_7__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__62_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__6_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__6_ccff_tail),
    .chany_top_out(sb_1__3__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__6_ccff_tail)
  );


  sb_1__3_
  sb_7__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__68_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__7_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__7_ccff_tail),
    .chany_top_out(sb_1__3__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__7_ccff_tail)
  );


  sb_1__3_
  sb_9__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__82_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__8_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__8_ccff_tail),
    .chany_top_out(sb_1__3__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__8_ccff_tail)
  );


  sb_1__3_
  sb_9__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__88_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__9_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__9_ccff_tail),
    .chany_top_out(sb_1__3__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__9_ccff_tail)
  );


  sb_1__3_
  sb_11__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__102_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__10_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__10_ccff_tail),
    .chany_top_out(sb_1__3__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__10_ccff_tail)
  );


  sb_1__3_
  sb_11__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__108_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__11_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__11_ccff_tail),
    .chany_top_out(sb_1__3__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__11_ccff_tail)
  );


  sb_1__12_
  sb_1__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__1_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__0_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_1_ccff_tail),
    .chanx_right_out(sb_1__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__0_ccff_tail)
  );


  sb_1__12_
  sb_2__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__2_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__1_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_2_ccff_tail),
    .chanx_right_out(sb_1__12__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__1_ccff_tail)
  );


  sb_1__12_
  sb_3__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__3_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__2_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_3_ccff_tail),
    .chanx_right_out(sb_1__12__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__2_ccff_tail)
  );


  sb_1__12_
  sb_4__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__4_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__3_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_4_ccff_tail),
    .chanx_right_out(sb_1__12__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__3_ccff_tail)
  );


  sb_1__12_
  sb_5__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__5_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__4_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_5_ccff_tail),
    .chanx_right_out(sb_1__12__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__4_ccff_tail)
  );


  sb_1__12_
  sb_6__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__6_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__59_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__5_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_6_ccff_tail),
    .chanx_right_out(sb_1__12__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__5_ccff_tail)
  );


  sb_1__12_
  sb_7__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__7_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__69_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__6_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_7_ccff_tail),
    .chanx_right_out(sb_1__12__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__6_ccff_tail)
  );


  sb_1__12_
  sb_8__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__8_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__79_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__7_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_8_ccff_tail),
    .chanx_right_out(sb_1__12__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__7_ccff_tail)
  );


  sb_1__12_
  sb_9__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__9_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__89_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__8_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_9_ccff_tail),
    .chanx_right_out(sb_1__12__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__8_ccff_tail)
  );


  sb_1__12_
  sb_10__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__10_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__99_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__9_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_10_ccff_tail),
    .chanx_right_out(sb_1__12__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__9_ccff_tail)
  );


  sb_1__12_
  sb_11__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_right_in(cbx_1__12__11_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__109_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__10_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_11_ccff_tail),
    .chanx_right_out(sb_1__12__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__10_ccff_tail)
  );


  sb_2__2_
  sb_2__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__10_ccff_tail),
    .chany_top_out(sb_2__2__0_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__0_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__0_ccff_tail)
  );


  sb_2__2_
  sb_2__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__16_ccff_tail),
    .chany_top_out(sb_2__2__1_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__1_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__1_ccff_tail)
  );


  sb_2__2_
  sb_4__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__28_ccff_tail),
    .chany_top_out(sb_2__2__2_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__2_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__2_ccff_tail)
  );


  sb_2__2_
  sb_4__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__34_ccff_tail),
    .chany_top_out(sb_2__2__3_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__3_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__3_ccff_tail)
  );


  sb_2__2_
  sb_6__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__46_ccff_tail),
    .chany_top_out(sb_2__2__4_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__4_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__4_ccff_tail)
  );


  sb_2__2_
  sb_6__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__61_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__57_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__52_ccff_tail),
    .chany_top_out(sb_2__2__5_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__5_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__5_ccff_tail)
  );


  sb_2__2_
  sb_8__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__73_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__71_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__64_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__64_ccff_tail),
    .chany_top_out(sb_2__2__6_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__6_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__6_ccff_tail)
  );


  sb_2__2_
  sb_8__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__79_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__77_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__70_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__70_ccff_tail),
    .chany_top_out(sb_2__2__7_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__7_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__7_ccff_tail)
  );


  sb_2__2_
  sb_10__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__91_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__91_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__82_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__82_ccff_tail),
    .chany_top_out(sb_2__2__8_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__8_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__8_ccff_tail)
  );


  sb_2__2_
  sb_10__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_2__3__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__97_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__97_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__88_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__88_ccff_tail),
    .chany_top_out(sb_2__2__9_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__9_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__9_ccff_tail)
  );


  sb_2__3_
  sb_2__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__0_ccff_tail),
    .chany_top_out(sb_2__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__0_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__0_ccff_tail)
  );


  sb_2__3_
  sb_2__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__1_ccff_tail),
    .chany_top_out(sb_2__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__1_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__1_ccff_tail)
  );


  sb_2__3_
  sb_4__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__2_ccff_tail),
    .chany_top_out(sb_2__3__2_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__2_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__2_ccff_tail)
  );


  sb_2__3_
  sb_4__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__3_ccff_tail),
    .chany_top_out(sb_2__3__3_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__3_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__3_ccff_tail)
  );


  sb_2__3_
  sb_6__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__4_ccff_tail),
    .chany_top_out(sb_2__3__4_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__4_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__4_ccff_tail)
  );


  sb_2__3_
  sb_6__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__58_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__5_ccff_tail),
    .chany_top_out(sb_2__3__5_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__5_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__5_ccff_tail)
  );


  sb_2__3_
  sb_8__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__72_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__6_ccff_tail),
    .chany_top_out(sb_2__3__6_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__6_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__6_ccff_tail)
  );


  sb_2__3_
  sb_8__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__78_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__7_ccff_tail),
    .chany_top_out(sb_2__3__7_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__7_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__7_ccff_tail)
  );


  sb_2__3_
  sb_10__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__92_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__8_ccff_tail),
    .chany_top_out(sb_2__3__8_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__8_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__8_ccff_tail)
  );


  sb_2__3_
  sb_10__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_1__1__98_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__9_ccff_tail),
    .chany_top_out(sb_2__3__9_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__9_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__9_ccff_tail)
  );


  sb_12__0_
  sb_12__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_left_in(cbx_1__0__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_0_ccff_tail),
    .chany_top_out(sb_12__0__0_chany_top_out[0:19]),
    .chanx_left_out(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[11])
  );


  sb_12__1_
  sb_12__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__0_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__99_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__99_ccff_tail),
    .chany_top_out(sb_12__1__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[10])
  );


  sb_12__1_
  sb_12__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__2_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__101_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__101_ccff_tail),
    .chany_top_out(sb_12__1__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[7])
  );


  sb_12__1_
  sb_12__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__3_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__102_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__102_ccff_tail),
    .chany_top_out(sb_12__1__2_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[6])
  );


  sb_12__1_
  sb_12__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__4_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__103_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__103_ccff_tail),
    .chany_top_out(sb_12__1__3_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[5])
  );


  sb_12__1_
  sb_12__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__5_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__104_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__104_ccff_tail),
    .chany_top_out(sb_12__1__4_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[4])
  );


  sb_12__1_
  sb_12__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__6_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__105_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__105_ccff_tail),
    .chany_top_out(sb_12__1__5_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[3])
  );


  sb_12__1_
  sb_12__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__8_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__107_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__107_ccff_tail),
    .chany_top_out(sb_12__1__6_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[0])
  );


  sb_12__2_
  sb_12__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__3__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__1_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__100_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__100_ccff_tail),
    .chany_top_out(sb_12__2__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__2__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[9])
  );


  sb_12__2_
  sb_12__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__3__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__7_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__106_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__106_ccff_tail),
    .chany_top_out(sb_12__2__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__2__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[2])
  );


  sb_12__3_
  sb_12__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__3__0_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__10_ccff_tail),
    .chany_top_out(sb_12__3__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__3__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[8])
  );


  sb_12__3_
  sb_12__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_top_in(cby_12__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__3__1_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__11_ccff_tail),
    .chany_top_out(sb_12__3__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__3__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[1])
  );


  sb_12__12_
  sb_12__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(cby_12__1__9_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__11_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(ccff_head[0]),
    .chany_bottom_out(sb_12__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_12__12__0_ccff_tail)
  );


  cbx_1__0_
  cbx_1__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__0__0_ccff_tail),
    .chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__0_ccff_tail)
  );


  cbx_1__0_
  cbx_2__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__0_ccff_tail),
    .chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__1_ccff_tail)
  );


  cbx_1__0_
  cbx_3__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__1_ccff_tail),
    .chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__2_ccff_tail)
  );


  cbx_1__0_
  cbx_4__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__2_ccff_tail),
    .chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__3_ccff_tail)
  );


  cbx_1__0_
  cbx_5__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__3_ccff_tail),
    .chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__4_ccff_tail)
  );


  cbx_1__0_
  cbx_6__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__4_ccff_tail),
    .chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__5_ccff_tail)
  );


  cbx_1__0_
  cbx_7__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__5_ccff_tail),
    .chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__6_ccff_tail)
  );


  cbx_1__0_
  cbx_8__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__6_ccff_tail),
    .chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__7_ccff_tail)
  );


  cbx_1__0_
  cbx_9__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__7_ccff_tail),
    .chanx_left_out(cbx_1__0__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__8_ccff_tail)
  );


  cbx_1__0_
  cbx_10__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__8_ccff_tail),
    .chanx_left_out(cbx_1__0__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__9_ccff_tail)
  );


  cbx_1__0_
  cbx_11__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__9_ccff_tail),
    .chanx_left_out(cbx_1__0__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__10_ccff_tail)
  );


  cbx_1__0_
  cbx_12__0_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__10_ccff_tail),
    .chanx_left_out(cbx_1__0__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
    .ccff_tail(cbx_1__0__11_ccff_tail)
  );


  cbx_1__1_
  cbx_1__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__0_ccff_tail),
    .chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__0_ccff_tail)
  );


  cbx_1__1_
  cbx_1__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__1_ccff_tail),
    .chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__1_ccff_tail)
  );


  cbx_1__1_
  cbx_1__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__2_ccff_tail),
    .chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__2_ccff_tail)
  );


  cbx_1__1_
  cbx_1__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__3_ccff_tail),
    .chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__3_ccff_tail)
  );


  cbx_1__1_
  cbx_1__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__4_ccff_tail),
    .chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__4_ccff_tail)
  );


  cbx_1__1_
  cbx_1__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__5_ccff_tail),
    .chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__5_ccff_tail)
  );


  cbx_1__1_
  cbx_1__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__6_ccff_tail),
    .chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__6_ccff_tail)
  );


  cbx_1__1_
  cbx_1__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__7_ccff_tail),
    .chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__7_ccff_tail)
  );


  cbx_1__1_
  cbx_1__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__8_ccff_tail),
    .chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__8_ccff_tail)
  );


  cbx_1__1_
  cbx_2__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__0_ccff_tail),
    .chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__9_ccff_tail)
  );


  cbx_1__1_
  cbx_2__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__0_ccff_tail),
    .chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__10_ccff_tail)
  );


  cbx_1__1_
  cbx_2__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__1_ccff_tail),
    .chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__11_ccff_tail)
  );


  cbx_1__1_
  cbx_2__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__2_ccff_tail),
    .chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__12_ccff_tail)
  );


  cbx_1__1_
  cbx_2__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__3_ccff_tail),
    .chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__13_ccff_tail)
  );


  cbx_1__1_
  cbx_2__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__4_ccff_tail),
    .chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__14_ccff_tail)
  );


  cbx_1__1_
  cbx_2__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__5_ccff_tail),
    .chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__15_ccff_tail)
  );


  cbx_1__1_
  cbx_2__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__1_ccff_tail),
    .chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__16_ccff_tail)
  );


  cbx_1__1_
  cbx_2__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__6_ccff_tail),
    .chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__17_ccff_tail)
  );


  cbx_1__1_
  cbx_3__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__7_ccff_tail),
    .chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__18_ccff_tail)
  );


  cbx_1__1_
  cbx_3__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__2_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__0_ccff_tail),
    .chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__19_ccff_tail)
  );


  cbx_1__1_
  cbx_3__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__8_ccff_tail),
    .chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__20_ccff_tail)
  );


  cbx_1__1_
  cbx_3__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__9_ccff_tail),
    .chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__21_ccff_tail)
  );


  cbx_1__1_
  cbx_3__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__10_ccff_tail),
    .chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__22_ccff_tail)
  );


  cbx_1__1_
  cbx_3__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__11_ccff_tail),
    .chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__23_ccff_tail)
  );


  cbx_1__1_
  cbx_3__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__12_ccff_tail),
    .chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__24_ccff_tail)
  );


  cbx_1__1_
  cbx_3__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__3_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__1_ccff_tail),
    .chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__25_ccff_tail)
  );


  cbx_1__1_
  cbx_3__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__13_ccff_tail),
    .chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__26_ccff_tail)
  );


  cbx_1__1_
  cbx_4__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__14_ccff_tail),
    .chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__27_ccff_tail)
  );


  cbx_1__1_
  cbx_4__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__2_ccff_tail),
    .chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__28_ccff_tail)
  );


  cbx_1__1_
  cbx_4__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__15_ccff_tail),
    .chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__29_ccff_tail)
  );


  cbx_1__1_
  cbx_4__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__16_ccff_tail),
    .chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__30_ccff_tail)
  );


  cbx_1__1_
  cbx_4__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__17_ccff_tail),
    .chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__31_ccff_tail)
  );


  cbx_1__1_
  cbx_4__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__18_ccff_tail),
    .chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__32_ccff_tail)
  );


  cbx_1__1_
  cbx_4__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__19_ccff_tail),
    .chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__33_ccff_tail)
  );


  cbx_1__1_
  cbx_4__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__3_ccff_tail),
    .chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__34_ccff_tail)
  );


  cbx_1__1_
  cbx_4__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__20_ccff_tail),
    .chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__35_ccff_tail)
  );


  cbx_1__1_
  cbx_5__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__21_ccff_tail),
    .chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__36_ccff_tail)
  );


  cbx_1__1_
  cbx_5__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__4_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__2_ccff_tail),
    .chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__37_ccff_tail)
  );


  cbx_1__1_
  cbx_5__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__22_ccff_tail),
    .chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__38_ccff_tail)
  );


  cbx_1__1_
  cbx_5__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__23_ccff_tail),
    .chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__39_ccff_tail)
  );


  cbx_1__1_
  cbx_5__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__24_ccff_tail),
    .chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__40_ccff_tail)
  );


  cbx_1__1_
  cbx_5__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__25_ccff_tail),
    .chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__41_ccff_tail)
  );


  cbx_1__1_
  cbx_5__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__26_ccff_tail),
    .chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__42_ccff_tail)
  );


  cbx_1__1_
  cbx_5__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__5_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__3_ccff_tail),
    .chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__43_ccff_tail)
  );


  cbx_1__1_
  cbx_5__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__27_ccff_tail),
    .chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__44_ccff_tail)
  );


  cbx_1__1_
  cbx_6__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__28_ccff_tail),
    .chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__45_ccff_tail)
  );


  cbx_1__1_
  cbx_6__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__4_ccff_tail),
    .chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__46_ccff_tail)
  );


  cbx_1__1_
  cbx_6__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__29_ccff_tail),
    .chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__47_ccff_tail)
  );


  cbx_1__1_
  cbx_6__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__30_ccff_tail),
    .chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__48_ccff_tail)
  );


  cbx_1__1_
  cbx_6__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__31_ccff_tail),
    .chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__49_ccff_tail)
  );


  cbx_1__1_
  cbx_6__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__32_ccff_tail),
    .chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__50_ccff_tail)
  );


  cbx_1__1_
  cbx_6__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__33_ccff_tail),
    .chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__51_ccff_tail)
  );


  cbx_1__1_
  cbx_6__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__5_ccff_tail),
    .chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__52_ccff_tail)
  );


  cbx_1__1_
  cbx_6__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__34_ccff_tail),
    .chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__53_ccff_tail)
  );


  cbx_1__1_
  cbx_7__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__35_ccff_tail),
    .chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__54_ccff_tail)
  );


  cbx_1__1_
  cbx_7__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__6_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__4_ccff_tail),
    .chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__55_ccff_tail)
  );


  cbx_1__1_
  cbx_7__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__36_ccff_tail),
    .chanx_left_out(cbx_1__1__56_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__56_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__56_ccff_tail)
  );


  cbx_1__1_
  cbx_7__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__37_ccff_tail),
    .chanx_left_out(cbx_1__1__57_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__57_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__57_ccff_tail)
  );


  cbx_1__1_
  cbx_7__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__38_ccff_tail),
    .chanx_left_out(cbx_1__1__58_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__58_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__58_ccff_tail)
  );


  cbx_1__1_
  cbx_7__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__39_ccff_tail),
    .chanx_left_out(cbx_1__1__59_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__59_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__59_ccff_tail)
  );


  cbx_1__1_
  cbx_7__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__40_ccff_tail),
    .chanx_left_out(cbx_1__1__60_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__60_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__60_ccff_tail)
  );


  cbx_1__1_
  cbx_7__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__7_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__5_ccff_tail),
    .chanx_left_out(cbx_1__1__61_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__61_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__61_ccff_tail)
  );


  cbx_1__1_
  cbx_7__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__41_ccff_tail),
    .chanx_left_out(cbx_1__1__62_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__62_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__62_ccff_tail)
  );


  cbx_1__1_
  cbx_8__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__42_ccff_tail),
    .chanx_left_out(cbx_1__1__63_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__63_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__63_ccff_tail)
  );


  cbx_1__1_
  cbx_8__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__6_ccff_tail),
    .chanx_left_out(cbx_1__1__64_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__64_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__64_ccff_tail)
  );


  cbx_1__1_
  cbx_8__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__43_ccff_tail),
    .chanx_left_out(cbx_1__1__65_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__65_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__65_ccff_tail)
  );


  cbx_1__1_
  cbx_8__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__44_ccff_tail),
    .chanx_left_out(cbx_1__1__66_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__66_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__66_ccff_tail)
  );


  cbx_1__1_
  cbx_8__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__45_ccff_tail),
    .chanx_left_out(cbx_1__1__67_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__67_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__67_ccff_tail)
  );


  cbx_1__1_
  cbx_8__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__46_ccff_tail),
    .chanx_left_out(cbx_1__1__68_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__68_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__68_ccff_tail)
  );


  cbx_1__1_
  cbx_8__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__47_ccff_tail),
    .chanx_left_out(cbx_1__1__69_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__69_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__69_ccff_tail)
  );


  cbx_1__1_
  cbx_8__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__7_ccff_tail),
    .chanx_left_out(cbx_1__1__70_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__70_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__70_ccff_tail)
  );


  cbx_1__1_
  cbx_8__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__48_ccff_tail),
    .chanx_left_out(cbx_1__1__71_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__71_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__71_ccff_tail)
  );


  cbx_1__1_
  cbx_9__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__49_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__49_ccff_tail),
    .chanx_left_out(cbx_1__1__72_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__72_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__72_ccff_tail)
  );


  cbx_1__1_
  cbx_9__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__8_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__6_ccff_tail),
    .chanx_left_out(cbx_1__1__73_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__73_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__73_ccff_tail)
  );


  cbx_1__1_
  cbx_9__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__50_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__50_ccff_tail),
    .chanx_left_out(cbx_1__1__74_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__74_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__74_ccff_tail)
  );


  cbx_1__1_
  cbx_9__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__51_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__51_ccff_tail),
    .chanx_left_out(cbx_1__1__75_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__75_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__75_ccff_tail)
  );


  cbx_1__1_
  cbx_9__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__52_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__52_ccff_tail),
    .chanx_left_out(cbx_1__1__76_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__76_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__76_ccff_tail)
  );


  cbx_1__1_
  cbx_9__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__53_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__53_ccff_tail),
    .chanx_left_out(cbx_1__1__77_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__77_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__77_ccff_tail)
  );


  cbx_1__1_
  cbx_9__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__54_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__54_ccff_tail),
    .chanx_left_out(cbx_1__1__78_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__78_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__78_ccff_tail)
  );


  cbx_1__1_
  cbx_9__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__9_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__7_ccff_tail),
    .chanx_left_out(cbx_1__1__79_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__79_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__79_ccff_tail)
  );


  cbx_1__1_
  cbx_9__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__55_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__55_ccff_tail),
    .chanx_left_out(cbx_1__1__80_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__80_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__80_ccff_tail)
  );


  cbx_1__1_
  cbx_10__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__56_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__56_ccff_tail),
    .chanx_left_out(cbx_1__1__81_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__81_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__81_ccff_tail)
  );


  cbx_1__1_
  cbx_10__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__8_ccff_tail),
    .chanx_left_out(cbx_1__1__82_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__82_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__82_ccff_tail)
  );


  cbx_1__1_
  cbx_10__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__57_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__57_ccff_tail),
    .chanx_left_out(cbx_1__1__83_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__83_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__83_ccff_tail)
  );


  cbx_1__1_
  cbx_10__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__58_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__58_ccff_tail),
    .chanx_left_out(cbx_1__1__84_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__84_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__84_ccff_tail)
  );


  cbx_1__1_
  cbx_10__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__59_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__59_ccff_tail),
    .chanx_left_out(cbx_1__1__85_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__85_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__85_ccff_tail)
  );


  cbx_1__1_
  cbx_10__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__60_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__60_ccff_tail),
    .chanx_left_out(cbx_1__1__86_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__86_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__86_ccff_tail)
  );


  cbx_1__1_
  cbx_10__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__61_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__61_ccff_tail),
    .chanx_left_out(cbx_1__1__87_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__87_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__87_ccff_tail)
  );


  cbx_1__1_
  cbx_10__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__9_ccff_tail),
    .chanx_left_out(cbx_1__1__88_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__88_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__88_ccff_tail)
  );


  cbx_1__1_
  cbx_10__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__62_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__62_ccff_tail),
    .chanx_left_out(cbx_1__1__89_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__89_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__89_ccff_tail)
  );


  cbx_1__1_
  cbx_11__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__63_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__63_ccff_tail),
    .chanx_left_out(cbx_1__1__90_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__90_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__90_ccff_tail)
  );


  cbx_1__1_
  cbx_11__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__10_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__8_ccff_tail),
    .chanx_left_out(cbx_1__1__91_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__91_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__91_ccff_tail)
  );


  cbx_1__1_
  cbx_11__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__64_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__64_ccff_tail),
    .chanx_left_out(cbx_1__1__92_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__92_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__92_ccff_tail)
  );


  cbx_1__1_
  cbx_11__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__65_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__65_ccff_tail),
    .chanx_left_out(cbx_1__1__93_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__93_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__93_ccff_tail)
  );


  cbx_1__1_
  cbx_11__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__66_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__66_ccff_tail),
    .chanx_left_out(cbx_1__1__94_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__94_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__94_ccff_tail)
  );


  cbx_1__1_
  cbx_11__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__67_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__67_ccff_tail),
    .chanx_left_out(cbx_1__1__95_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__95_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__95_ccff_tail)
  );


  cbx_1__1_
  cbx_11__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__68_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__68_ccff_tail),
    .chanx_left_out(cbx_1__1__96_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__96_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__96_ccff_tail)
  );


  cbx_1__1_
  cbx_11__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__2__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__11_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__9_ccff_tail),
    .chanx_left_out(cbx_1__1__97_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__97_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__97_ccff_tail)
  );


  cbx_1__1_
  cbx_11__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__69_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__69_ccff_tail),
    .chanx_left_out(cbx_1__1__98_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__98_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__98_ccff_tail)
  );


  cbx_1__1_
  cbx_12__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__70_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__70_ccff_tail),
    .chanx_left_out(cbx_1__1__99_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__99_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__99_ccff_tail)
  );


  cbx_1__1_
  cbx_12__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__10_ccff_tail),
    .chanx_left_out(cbx_1__1__100_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__100_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__100_ccff_tail)
  );


  cbx_1__1_
  cbx_12__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__71_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__71_ccff_tail),
    .chanx_left_out(cbx_1__1__101_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__101_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__101_ccff_tail)
  );


  cbx_1__1_
  cbx_12__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__72_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__72_ccff_tail),
    .chanx_left_out(cbx_1__1__102_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__102_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__102_ccff_tail)
  );


  cbx_1__1_
  cbx_12__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__73_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__73_ccff_tail),
    .chanx_left_out(cbx_1__1__103_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__103_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__103_ccff_tail)
  );


  cbx_1__1_
  cbx_12__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__74_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__74_ccff_tail),
    .chanx_left_out(cbx_1__1__104_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__104_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__104_ccff_tail)
  );


  cbx_1__1_
  cbx_12__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__75_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__75_ccff_tail),
    .chanx_left_out(cbx_1__1__105_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__105_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__105_ccff_tail)
  );


  cbx_1__1_
  cbx_12__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__2__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__11_ccff_tail),
    .chanx_left_out(cbx_1__1__106_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__106_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__106_ccff_tail)
  );


  cbx_1__1_
  cbx_12__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__1__76_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__76_ccff_tail),
    .chanx_left_out(cbx_1__1__107_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__107_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__107_ccff_tail)
  );


  cbx_1__3_
  cbx_1__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__3__0_ccff_tail),
    .chanx_left_out(cbx_1__3__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__0_ccff_tail)
  );


  cbx_1__3_
  cbx_1__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__3__1_ccff_tail),
    .chanx_left_out(cbx_1__3__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__1_ccff_tail)
  );


  cbx_1__3_
  cbx_3__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__2_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__0_ccff_tail),
    .chanx_left_out(cbx_1__3__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__2_ccff_tail)
  );


  cbx_1__3_
  cbx_3__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__3_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__1_ccff_tail),
    .chanx_left_out(cbx_1__3__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__3_ccff_tail)
  );


  cbx_1__3_
  cbx_5__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__4_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__2_ccff_tail),
    .chanx_left_out(cbx_1__3__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__4_ccff_tail)
  );


  cbx_1__3_
  cbx_5__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__5_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__3_ccff_tail),
    .chanx_left_out(cbx_1__3__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__5_ccff_tail)
  );


  cbx_1__3_
  cbx_7__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__6_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__4_ccff_tail),
    .chanx_left_out(cbx_1__3__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__6_ccff_tail)
  );


  cbx_1__3_
  cbx_7__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__7_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__5_ccff_tail),
    .chanx_left_out(cbx_1__3__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__7_ccff_tail)
  );


  cbx_1__3_
  cbx_9__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__8_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__6_ccff_tail),
    .chanx_left_out(cbx_1__3__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__8_ccff_tail)
  );


  cbx_1__3_
  cbx_9__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__9_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__7_ccff_tail),
    .chanx_left_out(cbx_1__3__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__9_ccff_tail)
  );


  cbx_1__3_
  cbx_11__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__10_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__8_ccff_tail),
    .chanx_left_out(cbx_1__3__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__10_ccff_tail)
  );


  cbx_1__3_
  cbx_11__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_2__3__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__11_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__9_ccff_tail),
    .chanx_left_out(cbx_1__3__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__11_ccff_tail)
  );


  cbx_1__12_
  cbx_1__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_0__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_head(grid_clb_9_ccff_tail),
    .chanx_left_out(cbx_1__12__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__0_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__0_ccff_tail)
  );


  cbx_1__12_
  cbx_2__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_head(grid_clb_19_ccff_tail),
    .chanx_left_out(cbx_1__12__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__1_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__1_ccff_tail)
  );


  cbx_1__12_
  cbx_3__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_head(grid_clb_29_ccff_tail),
    .chanx_left_out(cbx_1__12__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__2_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__2_ccff_tail)
  );


  cbx_1__12_
  cbx_4__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_head(grid_clb_39_ccff_tail),
    .chanx_left_out(cbx_1__12__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__3_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__3_ccff_tail)
  );


  cbx_1__12_
  cbx_5__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_head(grid_clb_49_ccff_tail),
    .chanx_left_out(cbx_1__12__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__4_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__4_ccff_tail)
  );


  cbx_1__12_
  cbx_6__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_head(grid_clb_59_ccff_tail),
    .chanx_left_out(cbx_1__12__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__5_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__5_ccff_tail)
  );


  cbx_1__12_
  cbx_7__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_head(grid_clb_69_ccff_tail),
    .chanx_left_out(cbx_1__12__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__6_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__6_ccff_tail)
  );


  cbx_1__12_
  cbx_8__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_head(grid_clb_79_ccff_tail),
    .chanx_left_out(cbx_1__12__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__7_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__7_ccff_tail)
  );


  cbx_1__12_
  cbx_9__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_head(grid_clb_89_ccff_tail),
    .chanx_left_out(cbx_1__12__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__8_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__8_ccff_tail)
  );


  cbx_1__12_
  cbx_10__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_head(grid_clb_99_ccff_tail),
    .chanx_left_out(cbx_1__12__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__9_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__9_ccff_tail)
  );


  cbx_1__12_
  cbx_11__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_head(grid_clb_109_ccff_tail),
    .chanx_left_out(cbx_1__12__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__10_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__10_ccff_tail)
  );


  cbx_1__12_
  cbx_12__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__12__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_head(grid_clb_119_ccff_tail),
    .chanx_left_out(cbx_1__12__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__11_chanx_right_out[0:19]),
    .top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__12__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__12__11_ccff_tail)
  );


  cbx_2__3_
  cbx_2__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__0_ccff_tail),
    .chanx_left_out(cbx_2__3__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__0_ccff_tail)
  );


  cbx_2__3_
  cbx_2__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__1_ccff_tail),
    .chanx_left_out(cbx_2__3__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__1_ccff_tail)
  );


  cbx_2__3_
  cbx_4__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__2_ccff_tail),
    .chanx_left_out(cbx_2__3__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__2_ccff_tail)
  );


  cbx_2__3_
  cbx_4__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__3_ccff_tail),
    .chanx_left_out(cbx_2__3__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__3_ccff_tail)
  );


  cbx_2__3_
  cbx_6__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__4_ccff_tail),
    .chanx_left_out(cbx_2__3__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__4_ccff_tail)
  );


  cbx_2__3_
  cbx_6__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__5_ccff_tail),
    .chanx_left_out(cbx_2__3__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__5_ccff_tail)
  );


  cbx_2__3_
  cbx_8__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__6_ccff_tail),
    .chanx_left_out(cbx_2__3__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__6_ccff_tail)
  );


  cbx_2__3_
  cbx_8__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__7_ccff_tail),
    .chanx_left_out(cbx_2__3__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__7_ccff_tail)
  );


  cbx_2__3_
  cbx_10__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__8_ccff_tail),
    .chanx_left_out(cbx_2__3__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__8_ccff_tail)
  );


  cbx_2__3_
  cbx_10__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__9_ccff_tail),
    .chanx_left_out(cbx_2__3__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__9_ccff_tail)
  );


  cbx_2__3_
  cbx_12__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__10_ccff_tail),
    .chanx_left_out(cbx_2__3__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__10_ccff_tail)
  );


  cbx_2__3_
  cbx_12__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chanx_left_in(sb_1__3__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__11_ccff_tail),
    .chanx_left_out(cbx_2__3__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__11_ccff_tail)
  );


  cby_0__1_
  cby_0__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_0_ccff_tail),
    .chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__0_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__0_ccff_tail)
  );


  cby_0__1_
  cby_0__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_1_ccff_tail),
    .chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__1_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__1_ccff_tail)
  );


  cby_0__1_
  cby_0__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__3__0_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_0_ccff_tail),
    .chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__2_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__2_ccff_tail)
  );


  cby_0__1_
  cby_0__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_2_ccff_tail),
    .chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__3_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__3_ccff_tail)
  );


  cby_0__1_
  cby_0__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_3_ccff_tail),
    .chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__4_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__4_ccff_tail)
  );


  cby_0__1_
  cby_0__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_4_ccff_tail),
    .chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__5_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__5_ccff_tail)
  );


  cby_0__1_
  cby_0__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_5_ccff_tail),
    .chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__6_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__6_ccff_tail)
  );


  cby_0__1_
  cby_0__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_6_ccff_tail),
    .chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__7_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__7_ccff_tail)
  );


  cby_0__1_
  cby_0__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_7_ccff_tail),
    .chany_bottom_out(cby_0__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__8_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__8_ccff_tail)
  );


  cby_0__1_
  cby_0__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_0__3__1_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_1_ccff_tail),
    .chany_bottom_out(cby_0__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__9_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__9_ccff_tail)
  );


  cby_0__1_
  cby_0__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_8_ccff_tail),
    .chany_bottom_out(cby_0__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__10_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__10_ccff_tail)
  );


  cby_0__1_
  cby_0__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_0__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__12__0_ccff_tail),
    .chany_bottom_out(cby_0__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__11_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
    .ccff_tail(cby_0__1__11_ccff_tail)
  );


  cby_1__1_
  cby_1__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_10_ccff_tail),
    .chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__0_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__0_ccff_tail)
  );


  cby_1__1_
  cby_1__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_11_ccff_tail),
    .chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__1_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__1_ccff_tail)
  );


  cby_1__1_
  cby_1__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_12_ccff_tail),
    .chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__2_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__2_ccff_tail)
  );


  cby_1__1_
  cby_1__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_13_ccff_tail),
    .chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__3_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__3_ccff_tail)
  );


  cby_1__1_
  cby_1__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_14_ccff_tail),
    .chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__4_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__4_ccff_tail)
  );


  cby_1__1_
  cby_1__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_15_ccff_tail),
    .chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__5_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__5_ccff_tail)
  );


  cby_1__1_
  cby_1__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_16_ccff_tail),
    .chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__6_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__6_ccff_tail)
  );


  cby_1__1_
  cby_1__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_17_ccff_tail),
    .chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__7_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__7_ccff_tail)
  );


  cby_1__1_
  cby_1__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_18_ccff_tail),
    .chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__8_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__8_ccff_tail)
  );


  cby_1__1_
  cby_1__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__0_ccff_tail),
    .chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__9_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__9_ccff_tail)
  );


  cby_1__1_
  cby_2__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_20_ccff_tail),
    .chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__10_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__10_ccff_tail)
  );


  cby_1__1_
  cby_2__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_21_ccff_tail),
    .chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__11_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__11_ccff_tail)
  );


  cby_1__1_
  cby_2__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_22_ccff_tail),
    .chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__12_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__12_ccff_tail)
  );


  cby_1__1_
  cby_2__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_23_ccff_tail),
    .chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__13_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__13_ccff_tail)
  );


  cby_1__1_
  cby_2__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_24_ccff_tail),
    .chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__14_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__14_ccff_tail)
  );


  cby_1__1_
  cby_2__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_25_ccff_tail),
    .chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__15_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__15_ccff_tail)
  );


  cby_1__1_
  cby_2__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_26_ccff_tail),
    .chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__16_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__16_ccff_tail)
  );


  cby_1__1_
  cby_2__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_27_ccff_tail),
    .chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__17_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__17_ccff_tail)
  );


  cby_1__1_
  cby_2__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_28_ccff_tail),
    .chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__18_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__18_ccff_tail)
  );


  cby_1__1_
  cby_2__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__1_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__1_ccff_tail),
    .chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__19_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__19_ccff_tail)
  );


  cby_1__1_
  cby_3__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_30_ccff_tail),
    .chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__20_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__20_ccff_tail)
  );


  cby_1__1_
  cby_3__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_31_ccff_tail),
    .chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__21_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__21_ccff_tail)
  );


  cby_1__1_
  cby_3__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_32_ccff_tail),
    .chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__22_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__22_ccff_tail)
  );


  cby_1__1_
  cby_3__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_33_ccff_tail),
    .chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__23_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__23_ccff_tail)
  );


  cby_1__1_
  cby_3__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_34_ccff_tail),
    .chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__24_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__24_ccff_tail)
  );


  cby_1__1_
  cby_3__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_35_ccff_tail),
    .chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__25_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__25_ccff_tail)
  );


  cby_1__1_
  cby_3__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_36_ccff_tail),
    .chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__26_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__26_ccff_tail)
  );


  cby_1__1_
  cby_3__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_37_ccff_tail),
    .chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__27_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__27_ccff_tail)
  );


  cby_1__1_
  cby_3__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_38_ccff_tail),
    .chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__28_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__28_ccff_tail)
  );


  cby_1__1_
  cby_3__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__2_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__2_ccff_tail),
    .chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__29_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__29_ccff_tail)
  );


  cby_1__1_
  cby_4__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_40_ccff_tail),
    .chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__30_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__30_ccff_tail)
  );


  cby_1__1_
  cby_4__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_41_ccff_tail),
    .chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__31_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__31_ccff_tail)
  );


  cby_1__1_
  cby_4__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_42_ccff_tail),
    .chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__32_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__32_ccff_tail)
  );


  cby_1__1_
  cby_4__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_43_ccff_tail),
    .chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__33_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__33_ccff_tail)
  );


  cby_1__1_
  cby_4__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_44_ccff_tail),
    .chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__34_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__34_ccff_tail)
  );


  cby_1__1_
  cby_4__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_45_ccff_tail),
    .chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__35_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__35_ccff_tail)
  );


  cby_1__1_
  cby_4__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_46_ccff_tail),
    .chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__36_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__36_ccff_tail)
  );


  cby_1__1_
  cby_4__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_47_ccff_tail),
    .chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__37_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__37_ccff_tail)
  );


  cby_1__1_
  cby_4__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_48_ccff_tail),
    .chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__38_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__38_ccff_tail)
  );


  cby_1__1_
  cby_4__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__3_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__3_ccff_tail),
    .chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__39_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__39_ccff_tail)
  );


  cby_1__1_
  cby_5__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_50_ccff_tail),
    .chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__40_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__40_ccff_tail)
  );


  cby_1__1_
  cby_5__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_51_ccff_tail),
    .chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__41_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__41_ccff_tail)
  );


  cby_1__1_
  cby_5__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_52_ccff_tail),
    .chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__42_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__42_ccff_tail)
  );


  cby_1__1_
  cby_5__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_53_ccff_tail),
    .chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__43_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__43_ccff_tail)
  );


  cby_1__1_
  cby_5__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_54_ccff_tail),
    .chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__44_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__44_ccff_tail)
  );


  cby_1__1_
  cby_5__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_55_ccff_tail),
    .chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__45_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__45_ccff_tail)
  );


  cby_1__1_
  cby_5__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_56_ccff_tail),
    .chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__46_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__46_ccff_tail)
  );


  cby_1__1_
  cby_5__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_57_ccff_tail),
    .chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__47_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__47_ccff_tail)
  );


  cby_1__1_
  cby_5__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_58_ccff_tail),
    .chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__48_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__48_ccff_tail)
  );


  cby_1__1_
  cby_5__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__4_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__4_ccff_tail),
    .chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__49_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__49_ccff_tail)
  );


  cby_1__1_
  cby_6__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_60_ccff_tail),
    .chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__50_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__50_ccff_tail)
  );


  cby_1__1_
  cby_6__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_61_ccff_tail),
    .chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__51_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__51_ccff_tail)
  );


  cby_1__1_
  cby_6__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_62_ccff_tail),
    .chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__52_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__52_ccff_tail)
  );


  cby_1__1_
  cby_6__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_63_ccff_tail),
    .chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__53_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__53_ccff_tail)
  );


  cby_1__1_
  cby_6__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_64_ccff_tail),
    .chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__54_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__54_ccff_tail)
  );


  cby_1__1_
  cby_6__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_65_ccff_tail),
    .chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__55_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__55_ccff_tail)
  );


  cby_1__1_
  cby_6__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_66_ccff_tail),
    .chany_bottom_out(cby_1__1__56_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__56_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__56_ccff_tail)
  );


  cby_1__1_
  cby_6__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_67_ccff_tail),
    .chany_bottom_out(cby_1__1__57_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__57_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__57_ccff_tail)
  );


  cby_1__1_
  cby_6__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_68_ccff_tail),
    .chany_bottom_out(cby_1__1__58_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__58_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__58_ccff_tail)
  );


  cby_1__1_
  cby_6__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__5_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__5_ccff_tail),
    .chany_bottom_out(cby_1__1__59_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__59_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__59_ccff_tail)
  );


  cby_1__1_
  cby_7__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_70_ccff_tail),
    .chany_bottom_out(cby_1__1__60_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__60_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__60_ccff_tail)
  );


  cby_1__1_
  cby_7__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_71_ccff_tail),
    .chany_bottom_out(cby_1__1__61_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__61_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__61_ccff_tail)
  );


  cby_1__1_
  cby_7__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_72_ccff_tail),
    .chany_bottom_out(cby_1__1__62_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__62_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__62_ccff_tail)
  );


  cby_1__1_
  cby_7__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_73_ccff_tail),
    .chany_bottom_out(cby_1__1__63_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__63_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__63_ccff_tail)
  );


  cby_1__1_
  cby_7__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_74_ccff_tail),
    .chany_bottom_out(cby_1__1__64_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__64_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__64_ccff_tail)
  );


  cby_1__1_
  cby_7__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_75_ccff_tail),
    .chany_bottom_out(cby_1__1__65_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__65_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__65_ccff_tail)
  );


  cby_1__1_
  cby_7__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_76_ccff_tail),
    .chany_bottom_out(cby_1__1__66_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__66_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__66_ccff_tail)
  );


  cby_1__1_
  cby_7__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_77_ccff_tail),
    .chany_bottom_out(cby_1__1__67_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__67_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__67_ccff_tail)
  );


  cby_1__1_
  cby_7__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_78_ccff_tail),
    .chany_bottom_out(cby_1__1__68_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__68_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__68_ccff_tail)
  );


  cby_1__1_
  cby_7__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__6_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__6_ccff_tail),
    .chany_bottom_out(cby_1__1__69_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__69_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__69_ccff_tail)
  );


  cby_1__1_
  cby_8__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__49_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_80_ccff_tail),
    .chany_bottom_out(cby_1__1__70_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__70_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__70_ccff_tail)
  );


  cby_1__1_
  cby_8__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__49_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_81_ccff_tail),
    .chany_bottom_out(cby_1__1__71_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__71_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__71_ccff_tail)
  );


  cby_1__1_
  cby_8__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__50_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_82_ccff_tail),
    .chany_bottom_out(cby_1__1__72_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__72_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__72_ccff_tail)
  );


  cby_1__1_
  cby_8__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__50_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__51_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_83_ccff_tail),
    .chany_bottom_out(cby_1__1__73_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__73_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__73_ccff_tail)
  );


  cby_1__1_
  cby_8__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__51_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__52_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_84_ccff_tail),
    .chany_bottom_out(cby_1__1__74_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__74_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__74_ccff_tail)
  );


  cby_1__1_
  cby_8__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__52_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__53_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_85_ccff_tail),
    .chany_bottom_out(cby_1__1__75_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__75_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__75_ccff_tail)
  );


  cby_1__1_
  cby_8__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__53_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__54_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_86_ccff_tail),
    .chany_bottom_out(cby_1__1__76_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__76_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__76_ccff_tail)
  );


  cby_1__1_
  cby_8__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__54_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_87_ccff_tail),
    .chany_bottom_out(cby_1__1__77_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__77_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__77_ccff_tail)
  );


  cby_1__1_
  cby_8__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__55_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_88_ccff_tail),
    .chany_bottom_out(cby_1__1__78_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__78_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__78_ccff_tail)
  );


  cby_1__1_
  cby_8__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__55_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__7_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__7_ccff_tail),
    .chany_bottom_out(cby_1__1__79_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__79_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__79_ccff_tail)
  );


  cby_1__1_
  cby_9__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__56_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_90_ccff_tail),
    .chany_bottom_out(cby_1__1__80_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__80_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__80_ccff_tail)
  );


  cby_1__1_
  cby_9__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__56_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_91_ccff_tail),
    .chany_bottom_out(cby_1__1__81_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__81_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__81_ccff_tail)
  );


  cby_1__1_
  cby_9__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__57_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_92_ccff_tail),
    .chany_bottom_out(cby_1__1__82_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__82_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__82_ccff_tail)
  );


  cby_1__1_
  cby_9__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__57_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__58_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_93_ccff_tail),
    .chany_bottom_out(cby_1__1__83_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__83_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__83_ccff_tail)
  );


  cby_1__1_
  cby_9__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__58_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__59_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_94_ccff_tail),
    .chany_bottom_out(cby_1__1__84_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__84_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__84_ccff_tail)
  );


  cby_1__1_
  cby_9__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__59_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__60_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_95_ccff_tail),
    .chany_bottom_out(cby_1__1__85_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__85_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__85_ccff_tail)
  );


  cby_1__1_
  cby_9__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__60_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__61_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_96_ccff_tail),
    .chany_bottom_out(cby_1__1__86_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__86_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__86_ccff_tail)
  );


  cby_1__1_
  cby_9__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__61_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_97_ccff_tail),
    .chany_bottom_out(cby_1__1__87_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__87_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__87_ccff_tail)
  );


  cby_1__1_
  cby_9__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__62_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_98_ccff_tail),
    .chany_bottom_out(cby_1__1__88_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__88_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__88_ccff_tail)
  );


  cby_1__1_
  cby_9__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__62_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__8_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__8_ccff_tail),
    .chany_bottom_out(cby_1__1__89_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__89_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__89_ccff_tail)
  );


  cby_1__1_
  cby_10__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__63_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_100_ccff_tail),
    .chany_bottom_out(cby_1__1__90_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__90_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__90_ccff_tail)
  );


  cby_1__1_
  cby_10__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__63_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_101_ccff_tail),
    .chany_bottom_out(cby_1__1__91_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__91_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__91_ccff_tail)
  );


  cby_1__1_
  cby_10__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__64_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_102_ccff_tail),
    .chany_bottom_out(cby_1__1__92_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__92_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__92_ccff_tail)
  );


  cby_1__1_
  cby_10__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__64_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__65_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_103_ccff_tail),
    .chany_bottom_out(cby_1__1__93_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__93_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__93_ccff_tail)
  );


  cby_1__1_
  cby_10__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__65_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__66_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_104_ccff_tail),
    .chany_bottom_out(cby_1__1__94_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__94_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__94_ccff_tail)
  );


  cby_1__1_
  cby_10__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__66_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__67_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_105_ccff_tail),
    .chany_bottom_out(cby_1__1__95_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__95_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__95_ccff_tail)
  );


  cby_1__1_
  cby_10__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__67_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__68_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_106_ccff_tail),
    .chany_bottom_out(cby_1__1__96_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__96_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__96_ccff_tail)
  );


  cby_1__1_
  cby_10__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__68_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_107_ccff_tail),
    .chany_bottom_out(cby_1__1__97_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__97_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__97_ccff_tail)
  );


  cby_1__1_
  cby_10__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__3__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__69_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_108_ccff_tail),
    .chany_bottom_out(cby_1__1__98_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__98_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__98_ccff_tail)
  );


  cby_1__1_
  cby_10__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__69_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__9_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__9_ccff_tail),
    .chany_bottom_out(cby_1__1__99_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__99_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__99_ccff_tail)
  );


  cby_1__1_
  cby_11__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__0__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__70_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_110_ccff_tail),
    .chany_bottom_out(cby_1__1__100_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__100_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__100_ccff_tail)
  );


  cby_1__1_
  cby_11__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__70_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_111_ccff_tail),
    .chany_bottom_out(cby_1__1__101_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__101_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__101_ccff_tail)
  );


  cby_1__1_
  cby_11__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__71_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_112_ccff_tail),
    .chany_bottom_out(cby_1__1__102_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__102_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__102_ccff_tail)
  );


  cby_1__1_
  cby_11__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__71_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__72_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_113_ccff_tail),
    .chany_bottom_out(cby_1__1__103_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__103_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__103_ccff_tail)
  );


  cby_1__1_
  cby_11__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__72_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__73_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_114_ccff_tail),
    .chany_bottom_out(cby_1__1__104_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__104_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__104_ccff_tail)
  );


  cby_1__1_
  cby_11__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__73_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__74_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_115_ccff_tail),
    .chany_bottom_out(cby_1__1__105_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__105_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__105_ccff_tail)
  );


  cby_1__1_
  cby_11__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__74_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__75_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_116_ccff_tail),
    .chany_bottom_out(cby_1__1__106_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__106_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__106_ccff_tail)
  );


  cby_1__1_
  cby_11__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__75_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_117_ccff_tail),
    .chany_bottom_out(cby_1__1__107_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__107_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__107_ccff_tail)
  );


  cby_1__1_
  cby_11__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__3__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__76_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_118_ccff_tail),
    .chany_bottom_out(cby_1__1__108_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__108_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__108_ccff_tail)
  );


  cby_1__1_
  cby_11__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_1__1__76_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__10_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__10_ccff_tail),
    .chany_bottom_out(cby_1__1__109_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__109_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__109_ccff_tail)
  );


  cby_1__3_
  cby_1__3_
  (
    .chany_bottom_in(sb_1__2__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__0_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__0_chany_top_out[0:19])
  );


  cby_1__3_
  cby_1__10_
  (
    .chany_bottom_in(sb_1__2__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__1_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__1_chany_top_out[0:19])
  );


  cby_1__3_
  cby_3__3_
  (
    .chany_bottom_in(sb_1__2__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__2_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__2_chany_top_out[0:19])
  );


  cby_1__3_
  cby_3__10_
  (
    .chany_bottom_in(sb_1__2__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__3_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__3_chany_top_out[0:19])
  );


  cby_1__3_
  cby_5__3_
  (
    .chany_bottom_in(sb_1__2__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__4_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__4_chany_top_out[0:19])
  );


  cby_1__3_
  cby_5__10_
  (
    .chany_bottom_in(sb_1__2__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__5_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__5_chany_top_out[0:19])
  );


  cby_1__3_
  cby_7__3_
  (
    .chany_bottom_in(sb_1__2__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__6_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__6_chany_top_out[0:19])
  );


  cby_1__3_
  cby_7__10_
  (
    .chany_bottom_in(sb_1__2__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__7_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__7_chany_top_out[0:19])
  );


  cby_1__3_
  cby_9__3_
  (
    .chany_bottom_in(sb_1__2__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__8_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__8_chany_top_out[0:19])
  );


  cby_1__3_
  cby_9__10_
  (
    .chany_bottom_in(sb_1__2__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__9_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__9_chany_top_out[0:19])
  );


  cby_1__3_
  cby_11__3_
  (
    .chany_bottom_in(sb_1__2__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__10_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__10_chany_top_out[0:19])
  );


  cby_1__3_
  cby_11__10_
  (
    .chany_bottom_in(sb_1__2__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__3__11_chany_bottom_out[0:19]),
    .chany_bottom_out(cby_1__3__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__3__11_chany_top_out[0:19])
  );


  cby_2__3_
  cby_2__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__0_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__0_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_2_ccff_tail),
    .chany_bottom_out(cby_2__3__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__0_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__0_ccff_tail)
  );


  cby_2__3_
  cby_2__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__1_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__1_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_3_ccff_tail),
    .chany_bottom_out(cby_2__3__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__1_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__1_ccff_tail)
  );


  cby_2__3_
  cby_4__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__2_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__2_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_4_ccff_tail),
    .chany_bottom_out(cby_2__3__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__2_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__2_ccff_tail)
  );


  cby_2__3_
  cby_4__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__3_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__3_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_5_ccff_tail),
    .chany_bottom_out(cby_2__3__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__3_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__3_ccff_tail)
  );


  cby_2__3_
  cby_6__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__4_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__4_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_6_ccff_tail),
    .chany_bottom_out(cby_2__3__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__4_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__4_ccff_tail)
  );


  cby_2__3_
  cby_6__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__5_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__5_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_7_ccff_tail),
    .chany_bottom_out(cby_2__3__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__5_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__5_ccff_tail)
  );


  cby_2__3_
  cby_8__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__6_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__6_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_8_ccff_tail),
    .chany_bottom_out(cby_2__3__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__6_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__6_ccff_tail)
  );


  cby_2__3_
  cby_8__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__7_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__7_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_9_ccff_tail),
    .chany_bottom_out(cby_2__3__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__7_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__7_ccff_tail)
  );


  cby_2__3_
  cby_10__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__8_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__8_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_10_ccff_tail),
    .chany_bottom_out(cby_2__3__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__8_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__8_ccff_tail)
  );


  cby_2__3_
  cby_10__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_2__2__9_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__9_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_11_ccff_tail),
    .chany_bottom_out(cby_2__3__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__9_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__9_ccff_tail)
  );


  cby_12__1_
  cby_12__1_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[11]),
    .chany_bottom_out(cby_12__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__0_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__0_ccff_tail)
  );


  cby_12__1_
  cby_12__2_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__2__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[10]),
    .chany_bottom_out(cby_12__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__1_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__1_ccff_tail)
  );


  cby_12__1_
  cby_12__4_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[8]),
    .chany_bottom_out(cby_12__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__2_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__2_ccff_tail)
  );


  cby_12__1_
  cby_12__5_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__2_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[7]),
    .chany_bottom_out(cby_12__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__3_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__3_ccff_tail)
  );


  cby_12__1_
  cby_12__6_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__3_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[6]),
    .chany_bottom_out(cby_12__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__4_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__4_ccff_tail)
  );


  cby_12__1_
  cby_12__7_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__4_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[5]),
    .chany_bottom_out(cby_12__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__5_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__5_ccff_tail)
  );


  cby_12__1_
  cby_12__8_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__5_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[4]),
    .chany_bottom_out(cby_12__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__6_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__6_ccff_tail)
  );


  cby_12__1_
  cby_12__9_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_12__2__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[3]),
    .chany_bottom_out(cby_12__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__7_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__7_ccff_tail)
  );


  cby_12__1_
  cby_12__11_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__6_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[1]),
    .chany_bottom_out(cby_12__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__8_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__8_ccff_tail)
  );


  cby_12__1_
  cby_12__12_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_12__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_12__12__0_ccff_tail),
    .chany_bottom_out(cby_12__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__9_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_12__1__9_ccff_tail)
  );


  cby_12__3_
  cby_12__3_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__2__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__3__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[9]),
    .chany_bottom_out(cby_12__3__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__3__0_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_12__3__0_ccff_tail)
  );


  cby_12__3_
  cby_12__10_
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .chany_bottom_in(sb_12__2__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__3__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[2]),
    .chany_bottom_out(cby_12__3__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__3__1_chany_top_out[0:19]),
    .right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_12__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_12__3__1_ccff_tail)
  );


  direct_interc
  direct_interc_0_
  (
    .in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_0_out)
  );


  direct_interc
  direct_interc_1_
  (
    .in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_1_out)
  );


  direct_interc
  direct_interc_2_
  (
    .in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_2_out)
  );


  direct_interc
  direct_interc_3_
  (
    .in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_3_out)
  );


  direct_interc
  direct_interc_4_
  (
    .in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_4_out)
  );


  direct_interc
  direct_interc_5_
  (
    .in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_5_out)
  );


  direct_interc
  direct_interc_6_
  (
    .in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_6_out)
  );


  direct_interc
  direct_interc_7_
  (
    .in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_7_out)
  );


  direct_interc
  direct_interc_8_
  (
    .in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_8_out)
  );


  direct_interc
  direct_interc_9_
  (
    .in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_9_out)
  );


  direct_interc
  direct_interc_10_
  (
    .in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_10_out)
  );


  direct_interc
  direct_interc_11_
  (
    .in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_11_out)
  );


  direct_interc
  direct_interc_12_
  (
    .in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_12_out)
  );


  direct_interc
  direct_interc_13_
  (
    .in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_13_out)
  );


  direct_interc
  direct_interc_14_
  (
    .in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_14_out)
  );


  direct_interc
  direct_interc_15_
  (
    .in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_15_out)
  );


  direct_interc
  direct_interc_16_
  (
    .in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_16_out)
  );


  direct_interc
  direct_interc_17_
  (
    .in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_17_out)
  );


  direct_interc
  direct_interc_18_
  (
    .in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_18_out)
  );


  direct_interc
  direct_interc_19_
  (
    .in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_19_out)
  );


  direct_interc
  direct_interc_20_
  (
    .in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_20_out)
  );


  direct_interc
  direct_interc_21_
  (
    .in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_21_out)
  );


  direct_interc
  direct_interc_22_
  (
    .in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_22_out)
  );


  direct_interc
  direct_interc_23_
  (
    .in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_23_out)
  );


  direct_interc
  direct_interc_24_
  (
    .in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_24_out)
  );


  direct_interc
  direct_interc_25_
  (
    .in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_25_out)
  );


  direct_interc
  direct_interc_26_
  (
    .in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_26_out)
  );


  direct_interc
  direct_interc_27_
  (
    .in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_27_out)
  );


  direct_interc
  direct_interc_28_
  (
    .in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_28_out)
  );


  direct_interc
  direct_interc_29_
  (
    .in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_29_out)
  );


  direct_interc
  direct_interc_30_
  (
    .in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_30_out)
  );


  direct_interc
  direct_interc_31_
  (
    .in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_31_out)
  );


  direct_interc
  direct_interc_32_
  (
    .in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_32_out)
  );


  direct_interc
  direct_interc_33_
  (
    .in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_33_out)
  );


  direct_interc
  direct_interc_34_
  (
    .in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_34_out)
  );


  direct_interc
  direct_interc_35_
  (
    .in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_35_out)
  );


  direct_interc
  direct_interc_36_
  (
    .in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_36_out)
  );


  direct_interc
  direct_interc_37_
  (
    .in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_37_out)
  );


  direct_interc
  direct_interc_38_
  (
    .in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_38_out)
  );


  direct_interc
  direct_interc_39_
  (
    .in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_39_out)
  );


  direct_interc
  direct_interc_40_
  (
    .in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_40_out)
  );


  direct_interc
  direct_interc_41_
  (
    .in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_41_out)
  );


  direct_interc
  direct_interc_42_
  (
    .in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_42_out)
  );


  direct_interc
  direct_interc_43_
  (
    .in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_43_out)
  );


  direct_interc
  direct_interc_44_
  (
    .in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_44_out)
  );


  direct_interc
  direct_interc_45_
  (
    .in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_45_out)
  );


  direct_interc
  direct_interc_46_
  (
    .in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_46_out)
  );


  direct_interc
  direct_interc_47_
  (
    .in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_47_out)
  );


  direct_interc
  direct_interc_48_
  (
    .in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_48_out)
  );


  direct_interc
  direct_interc_49_
  (
    .in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_49_out)
  );


  direct_interc
  direct_interc_50_
  (
    .in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_50_out)
  );


  direct_interc
  direct_interc_51_
  (
    .in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_51_out)
  );


  direct_interc
  direct_interc_52_
  (
    .in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_52_out)
  );


  direct_interc
  direct_interc_53_
  (
    .in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_53_out)
  );


  direct_interc
  direct_interc_54_
  (
    .in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_54_out)
  );


  direct_interc
  direct_interc_55_
  (
    .in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_55_out)
  );


  direct_interc
  direct_interc_56_
  (
    .in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_56_out)
  );


  direct_interc
  direct_interc_57_
  (
    .in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_57_out)
  );


  direct_interc
  direct_interc_58_
  (
    .in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_58_out)
  );


  direct_interc
  direct_interc_59_
  (
    .in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_59_out)
  );


  direct_interc
  direct_interc_60_
  (
    .in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_60_out)
  );


  direct_interc
  direct_interc_61_
  (
    .in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_61_out)
  );


  direct_interc
  direct_interc_62_
  (
    .in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_62_out)
  );


  direct_interc
  direct_interc_63_
  (
    .in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_63_out)
  );


  direct_interc
  direct_interc_64_
  (
    .in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_64_out)
  );


  direct_interc
  direct_interc_65_
  (
    .in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_65_out)
  );


  direct_interc
  direct_interc_66_
  (
    .in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_66_out)
  );


  direct_interc
  direct_interc_67_
  (
    .in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_67_out)
  );


  direct_interc
  direct_interc_68_
  (
    .in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_68_out)
  );


  direct_interc
  direct_interc_69_
  (
    .in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_69_out)
  );


  direct_interc
  direct_interc_70_
  (
    .in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_70_out)
  );


  direct_interc
  direct_interc_71_
  (
    .in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_71_out)
  );


  direct_interc
  direct_interc_72_
  (
    .in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_72_out)
  );


  direct_interc
  direct_interc_73_
  (
    .in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_73_out)
  );


  direct_interc
  direct_interc_74_
  (
    .in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_74_out)
  );


  direct_interc
  direct_interc_75_
  (
    .in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_75_out)
  );


  direct_interc
  direct_interc_76_
  (
    .in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_76_out)
  );


  direct_interc
  direct_interc_77_
  (
    .in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_77_out)
  );


  direct_interc
  direct_interc_78_
  (
    .in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_78_out)
  );


  direct_interc
  direct_interc_79_
  (
    .in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_79_out)
  );


  direct_interc
  direct_interc_80_
  (
    .in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_80_out)
  );


  direct_interc
  direct_interc_81_
  (
    .in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_81_out)
  );


  direct_interc
  direct_interc_82_
  (
    .in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_82_out)
  );


  direct_interc
  direct_interc_83_
  (
    .in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_83_out)
  );


  direct_interc
  direct_interc_84_
  (
    .in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_84_out)
  );


  direct_interc
  direct_interc_85_
  (
    .in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_85_out)
  );


  direct_interc
  direct_interc_86_
  (
    .in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_86_out)
  );


  direct_interc
  direct_interc_87_
  (
    .in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_87_out)
  );


  direct_interc
  direct_interc_88_
  (
    .in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_88_out)
  );


  direct_interc
  direct_interc_89_
  (
    .in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_89_out)
  );


  direct_interc
  direct_interc_90_
  (
    .in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_90_out)
  );


  direct_interc
  direct_interc_91_
  (
    .in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_91_out)
  );


  direct_interc
  direct_interc_92_
  (
    .in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_92_out)
  );


  direct_interc
  direct_interc_93_
  (
    .in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_93_out)
  );


  direct_interc
  direct_interc_94_
  (
    .in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_94_out)
  );


  direct_interc
  direct_interc_95_
  (
    .in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_95_out)
  );


  direct_interc
  direct_interc_96_
  (
    .in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_96_out)
  );


  direct_interc
  direct_interc_97_
  (
    .in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_97_out)
  );


  direct_interc
  direct_interc_98_
  (
    .in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_98_out)
  );


  direct_interc
  direct_interc_99_
  (
    .in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_99_out)
  );


  direct_interc
  direct_interc_100_
  (
    .in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_100_out)
  );


  direct_interc
  direct_interc_101_
  (
    .in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_101_out)
  );


  direct_interc
  direct_interc_102_
  (
    .in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_102_out)
  );


  direct_interc
  direct_interc_103_
  (
    .in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_103_out)
  );


  direct_interc
  direct_interc_104_
  (
    .in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_104_out)
  );


  direct_interc
  direct_interc_105_
  (
    .in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_105_out)
  );


  direct_interc
  direct_interc_106_
  (
    .in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_106_out)
  );


  direct_interc
  direct_interc_107_
  (
    .in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_107_out)
  );


  direct_interc
  direct_interc_108_
  (
    .in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_108_out)
  );


  direct_interc
  direct_interc_109_
  (
    .in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_109_out)
  );


  direct_interc
  direct_interc_110_
  (
    .in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_110_out)
  );


  direct_interc
  direct_interc_111_
  (
    .in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_111_out)
  );


  direct_interc
  direct_interc_112_
  (
    .in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_112_out)
  );


  direct_interc
  direct_interc_113_
  (
    .in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_113_out)
  );


  direct_interc
  direct_interc_114_
  (
    .in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_114_out)
  );


  direct_interc
  direct_interc_115_
  (
    .in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_115_out)
  );


  direct_interc
  direct_interc_116_
  (
    .in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_116_out)
  );


  direct_interc
  direct_interc_117_
  (
    .in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_117_out)
  );


  direct_interc
  direct_interc_118_
  (
    .in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_118_out)
  );


  direct_interc
  direct_interc_119_
  (
    .in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_119_out)
  );


  direct_interc
  direct_interc_120_
  (
    .in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_120_out)
  );


  direct_interc
  direct_interc_121_
  (
    .in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_121_out)
  );


  direct_interc
  direct_interc_122_
  (
    .in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_122_out)
  );


  direct_interc
  direct_interc_123_
  (
    .in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_123_out)
  );


  direct_interc
  direct_interc_124_
  (
    .in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_124_out)
  );


  direct_interc
  direct_interc_125_
  (
    .in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_125_out)
  );


  direct_interc
  direct_interc_126_
  (
    .in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_126_out)
  );


  direct_interc
  direct_interc_127_
  (
    .in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_127_out)
  );


  direct_interc
  direct_interc_128_
  (
    .in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_128_out)
  );


  direct_interc
  direct_interc_129_
  (
    .in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_129_out)
  );


  direct_interc
  direct_interc_130_
  (
    .in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_130_out)
  );


  direct_interc
  direct_interc_131_
  (
    .in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_131_out)
  );


  direct_interc
  direct_interc_132_
  (
    .in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_132_out)
  );


  direct_interc
  direct_interc_133_
  (
    .in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_133_out)
  );


  direct_interc
  direct_interc_134_
  (
    .in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_134_out)
  );


  direct_interc
  direct_interc_135_
  (
    .in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_135_out)
  );


  direct_interc
  direct_interc_136_
  (
    .in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_136_out)
  );


  direct_interc
  direct_interc_137_
  (
    .in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_137_out)
  );


  direct_interc
  direct_interc_138_
  (
    .in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_138_out)
  );


  direct_interc
  direct_interc_139_
  (
    .in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_139_out)
  );


  direct_interc
  direct_interc_140_
  (
    .in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_140_out)
  );


  direct_interc
  direct_interc_141_
  (
    .in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_141_out)
  );


  direct_interc
  direct_interc_142_
  (
    .in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_142_out)
  );


  direct_interc
  direct_interc_143_
  (
    .in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_143_out)
  );


  direct_interc
  direct_interc_144_
  (
    .in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_144_out)
  );


  direct_interc
  direct_interc_145_
  (
    .in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_145_out)
  );


  direct_interc
  direct_interc_146_
  (
    .in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_146_out)
  );


  direct_interc
  direct_interc_147_
  (
    .in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_147_out)
  );


  direct_interc
  direct_interc_148_
  (
    .in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_148_out)
  );


  direct_interc
  direct_interc_149_
  (
    .in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_149_out)
  );


  direct_interc
  direct_interc_150_
  (
    .in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_150_out)
  );


  direct_interc
  direct_interc_151_
  (
    .in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_151_out)
  );


  direct_interc
  direct_interc_152_
  (
    .in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_152_out)
  );


  direct_interc
  direct_interc_153_
  (
    .in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_153_out)
  );


  direct_interc
  direct_interc_154_
  (
    .in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_154_out)
  );


  direct_interc
  direct_interc_155_
  (
    .in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_155_out)
  );


  direct_interc
  direct_interc_156_
  (
    .in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_156_out)
  );


  direct_interc
  direct_interc_157_
  (
    .in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_157_out)
  );


  direct_interc
  direct_interc_158_
  (
    .in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_158_out)
  );


  direct_interc
  direct_interc_159_
  (
    .in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_159_out)
  );


  direct_interc
  direct_interc_160_
  (
    .in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_160_out)
  );


  direct_interc
  direct_interc_161_
  (
    .in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_161_out)
  );


  direct_interc
  direct_interc_162_
  (
    .in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_162_out)
  );


  direct_interc
  direct_interc_163_
  (
    .in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_163_out)
  );


  direct_interc
  direct_interc_164_
  (
    .in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_164_out)
  );


  direct_interc
  direct_interc_165_
  (
    .in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_165_out)
  );


  direct_interc
  direct_interc_166_
  (
    .in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_166_out)
  );


  direct_interc
  direct_interc_167_
  (
    .in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_167_out)
  );


  direct_interc
  direct_interc_168_
  (
    .in(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_168_out)
  );


  direct_interc
  direct_interc_169_
  (
    .in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_169_out)
  );


  direct_interc
  direct_interc_170_
  (
    .in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_170_out)
  );


  direct_interc
  direct_interc_171_
  (
    .in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_171_out)
  );


  direct_interc
  direct_interc_172_
  (
    .in(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_172_out)
  );


  direct_interc
  direct_interc_173_
  (
    .in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_173_out)
  );


  direct_interc
  direct_interc_174_
  (
    .in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_174_out)
  );


  direct_interc
  direct_interc_175_
  (
    .in(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_175_out)
  );


  direct_interc
  direct_interc_176_
  (
    .in(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_176_out)
  );


  direct_interc
  direct_interc_177_
  (
    .in(grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_177_out)
  );


  direct_interc
  direct_interc_178_
  (
    .in(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_178_out)
  );


endmodule

