//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
// `default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(config_enable,
                pReset,
                prog_clk,
                Test_en,
                IO_ISOL_N,
                clk,
                reset,
                gfpga_pad_sofa_plus_io_SOC_IN,
                gfpga_pad_sofa_plus_io_SOC_OUT,
                gfpga_pad_sofa_plus_io_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GPIN PORTS -----
input [0:175] gfpga_pad_sofa_plus_io_SOC_IN;
//----- GPOUT PORTS -----
output [0:175] gfpga_pad_sofa_plus_io_SOC_OUT;
//----- GPOUT PORTS -----
output [0:175] gfpga_pad_sofa_plus_io_SOC_DIR;
//----- INPUT PORTS -----
input [0:11] ccff_head;
//----- OUTPUT PORTS -----
output [0:11] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:63] cbx_1__0__0_chanx_left_out;
wire [0:63] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__100_ccff_tail;
wire [0:63] cbx_1__0__100_chanx_left_out;
wire [0:63] cbx_1__0__100_chanx_right_out;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__101_ccff_tail;
wire [0:63] cbx_1__0__101_chanx_left_out;
wire [0:63] cbx_1__0__101_chanx_right_out;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__102_ccff_tail;
wire [0:63] cbx_1__0__102_chanx_left_out;
wire [0:63] cbx_1__0__102_chanx_right_out;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__103_ccff_tail;
wire [0:63] cbx_1__0__103_chanx_left_out;
wire [0:63] cbx_1__0__103_chanx_right_out;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:63] cbx_1__0__104_chanx_left_out;
wire [0:63] cbx_1__0__104_chanx_right_out;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__105_ccff_tail;
wire [0:63] cbx_1__0__105_chanx_left_out;
wire [0:63] cbx_1__0__105_chanx_right_out;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__106_ccff_tail;
wire [0:63] cbx_1__0__106_chanx_left_out;
wire [0:63] cbx_1__0__106_chanx_right_out;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__107_ccff_tail;
wire [0:63] cbx_1__0__107_chanx_left_out;
wire [0:63] cbx_1__0__107_chanx_right_out;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__108_ccff_tail;
wire [0:63] cbx_1__0__108_chanx_left_out;
wire [0:63] cbx_1__0__108_chanx_right_out;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__109_ccff_tail;
wire [0:63] cbx_1__0__109_chanx_left_out;
wire [0:63] cbx_1__0__109_chanx_right_out;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__10_ccff_tail;
wire [0:63] cbx_1__0__10_chanx_left_out;
wire [0:63] cbx_1__0__10_chanx_right_out;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__110_ccff_tail;
wire [0:63] cbx_1__0__110_chanx_left_out;
wire [0:63] cbx_1__0__110_chanx_right_out;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__111_ccff_tail;
wire [0:63] cbx_1__0__111_chanx_left_out;
wire [0:63] cbx_1__0__111_chanx_right_out;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__112_ccff_tail;
wire [0:63] cbx_1__0__112_chanx_left_out;
wire [0:63] cbx_1__0__112_chanx_right_out;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__113_ccff_tail;
wire [0:63] cbx_1__0__113_chanx_left_out;
wire [0:63] cbx_1__0__113_chanx_right_out;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__114_ccff_tail;
wire [0:63] cbx_1__0__114_chanx_left_out;
wire [0:63] cbx_1__0__114_chanx_right_out;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__115_ccff_tail;
wire [0:63] cbx_1__0__115_chanx_left_out;
wire [0:63] cbx_1__0__115_chanx_right_out;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__116_ccff_tail;
wire [0:63] cbx_1__0__116_chanx_left_out;
wire [0:63] cbx_1__0__116_chanx_right_out;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__117_ccff_tail;
wire [0:63] cbx_1__0__117_chanx_left_out;
wire [0:63] cbx_1__0__117_chanx_right_out;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__118_ccff_tail;
wire [0:63] cbx_1__0__118_chanx_left_out;
wire [0:63] cbx_1__0__118_chanx_right_out;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__119_ccff_tail;
wire [0:63] cbx_1__0__119_chanx_left_out;
wire [0:63] cbx_1__0__119_chanx_right_out;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__11_ccff_tail;
wire [0:63] cbx_1__0__11_chanx_left_out;
wire [0:63] cbx_1__0__11_chanx_right_out;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__120_ccff_tail;
wire [0:63] cbx_1__0__120_chanx_left_out;
wire [0:63] cbx_1__0__120_chanx_right_out;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__121_ccff_tail;
wire [0:63] cbx_1__0__121_chanx_left_out;
wire [0:63] cbx_1__0__121_chanx_right_out;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__122_ccff_tail;
wire [0:63] cbx_1__0__122_chanx_left_out;
wire [0:63] cbx_1__0__122_chanx_right_out;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__123_ccff_tail;
wire [0:63] cbx_1__0__123_chanx_left_out;
wire [0:63] cbx_1__0__123_chanx_right_out;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__124_ccff_tail;
wire [0:63] cbx_1__0__124_chanx_left_out;
wire [0:63] cbx_1__0__124_chanx_right_out;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__125_ccff_tail;
wire [0:63] cbx_1__0__125_chanx_left_out;
wire [0:63] cbx_1__0__125_chanx_right_out;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__126_ccff_tail;
wire [0:63] cbx_1__0__126_chanx_left_out;
wire [0:63] cbx_1__0__126_chanx_right_out;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__127_ccff_tail;
wire [0:63] cbx_1__0__127_chanx_left_out;
wire [0:63] cbx_1__0__127_chanx_right_out;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__128_ccff_tail;
wire [0:63] cbx_1__0__128_chanx_left_out;
wire [0:63] cbx_1__0__128_chanx_right_out;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__129_ccff_tail;
wire [0:63] cbx_1__0__129_chanx_left_out;
wire [0:63] cbx_1__0__129_chanx_right_out;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__12_ccff_tail;
wire [0:63] cbx_1__0__12_chanx_left_out;
wire [0:63] cbx_1__0__12_chanx_right_out;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__130_ccff_tail;
wire [0:63] cbx_1__0__130_chanx_left_out;
wire [0:63] cbx_1__0__130_chanx_right_out;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__131_ccff_tail;
wire [0:63] cbx_1__0__131_chanx_left_out;
wire [0:63] cbx_1__0__131_chanx_right_out;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__132_ccff_tail;
wire [0:63] cbx_1__0__132_chanx_left_out;
wire [0:63] cbx_1__0__132_chanx_right_out;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__133_ccff_tail;
wire [0:63] cbx_1__0__133_chanx_left_out;
wire [0:63] cbx_1__0__133_chanx_right_out;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__134_ccff_tail;
wire [0:63] cbx_1__0__134_chanx_left_out;
wire [0:63] cbx_1__0__134_chanx_right_out;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__135_ccff_tail;
wire [0:63] cbx_1__0__135_chanx_left_out;
wire [0:63] cbx_1__0__135_chanx_right_out;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__136_ccff_tail;
wire [0:63] cbx_1__0__136_chanx_left_out;
wire [0:63] cbx_1__0__136_chanx_right_out;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__137_ccff_tail;
wire [0:63] cbx_1__0__137_chanx_left_out;
wire [0:63] cbx_1__0__137_chanx_right_out;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__138_ccff_tail;
wire [0:63] cbx_1__0__138_chanx_left_out;
wire [0:63] cbx_1__0__138_chanx_right_out;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__139_ccff_tail;
wire [0:63] cbx_1__0__139_chanx_left_out;
wire [0:63] cbx_1__0__139_chanx_right_out;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__13_ccff_tail;
wire [0:63] cbx_1__0__13_chanx_left_out;
wire [0:63] cbx_1__0__13_chanx_right_out;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__140_ccff_tail;
wire [0:63] cbx_1__0__140_chanx_left_out;
wire [0:63] cbx_1__0__140_chanx_right_out;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__141_ccff_tail;
wire [0:63] cbx_1__0__141_chanx_left_out;
wire [0:63] cbx_1__0__141_chanx_right_out;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__142_ccff_tail;
wire [0:63] cbx_1__0__142_chanx_left_out;
wire [0:63] cbx_1__0__142_chanx_right_out;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__143_ccff_tail;
wire [0:63] cbx_1__0__143_chanx_left_out;
wire [0:63] cbx_1__0__143_chanx_right_out;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__144_ccff_tail;
wire [0:63] cbx_1__0__144_chanx_left_out;
wire [0:63] cbx_1__0__144_chanx_right_out;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__145_ccff_tail;
wire [0:63] cbx_1__0__145_chanx_left_out;
wire [0:63] cbx_1__0__145_chanx_right_out;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__146_ccff_tail;
wire [0:63] cbx_1__0__146_chanx_left_out;
wire [0:63] cbx_1__0__146_chanx_right_out;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__147_ccff_tail;
wire [0:63] cbx_1__0__147_chanx_left_out;
wire [0:63] cbx_1__0__147_chanx_right_out;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__148_ccff_tail;
wire [0:63] cbx_1__0__148_chanx_left_out;
wire [0:63] cbx_1__0__148_chanx_right_out;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__149_ccff_tail;
wire [0:63] cbx_1__0__149_chanx_left_out;
wire [0:63] cbx_1__0__149_chanx_right_out;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__14_ccff_tail;
wire [0:63] cbx_1__0__14_chanx_left_out;
wire [0:63] cbx_1__0__14_chanx_right_out;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__150_ccff_tail;
wire [0:63] cbx_1__0__150_chanx_left_out;
wire [0:63] cbx_1__0__150_chanx_right_out;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__151_ccff_tail;
wire [0:63] cbx_1__0__151_chanx_left_out;
wire [0:63] cbx_1__0__151_chanx_right_out;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__152_ccff_tail;
wire [0:63] cbx_1__0__152_chanx_left_out;
wire [0:63] cbx_1__0__152_chanx_right_out;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__153_ccff_tail;
wire [0:63] cbx_1__0__153_chanx_left_out;
wire [0:63] cbx_1__0__153_chanx_right_out;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__154_ccff_tail;
wire [0:63] cbx_1__0__154_chanx_left_out;
wire [0:63] cbx_1__0__154_chanx_right_out;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__155_ccff_tail;
wire [0:63] cbx_1__0__155_chanx_left_out;
wire [0:63] cbx_1__0__155_chanx_right_out;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__156_ccff_tail;
wire [0:63] cbx_1__0__156_chanx_left_out;
wire [0:63] cbx_1__0__156_chanx_right_out;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__157_ccff_tail;
wire [0:63] cbx_1__0__157_chanx_left_out;
wire [0:63] cbx_1__0__157_chanx_right_out;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__158_ccff_tail;
wire [0:63] cbx_1__0__158_chanx_left_out;
wire [0:63] cbx_1__0__158_chanx_right_out;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__159_ccff_tail;
wire [0:63] cbx_1__0__159_chanx_left_out;
wire [0:63] cbx_1__0__159_chanx_right_out;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__15_ccff_tail;
wire [0:63] cbx_1__0__15_chanx_left_out;
wire [0:63] cbx_1__0__15_chanx_right_out;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__160_ccff_tail;
wire [0:63] cbx_1__0__160_chanx_left_out;
wire [0:63] cbx_1__0__160_chanx_right_out;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__161_ccff_tail;
wire [0:63] cbx_1__0__161_chanx_left_out;
wire [0:63] cbx_1__0__161_chanx_right_out;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__162_ccff_tail;
wire [0:63] cbx_1__0__162_chanx_left_out;
wire [0:63] cbx_1__0__162_chanx_right_out;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__163_ccff_tail;
wire [0:63] cbx_1__0__163_chanx_left_out;
wire [0:63] cbx_1__0__163_chanx_right_out;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__164_ccff_tail;
wire [0:63] cbx_1__0__164_chanx_left_out;
wire [0:63] cbx_1__0__164_chanx_right_out;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__165_ccff_tail;
wire [0:63] cbx_1__0__165_chanx_left_out;
wire [0:63] cbx_1__0__165_chanx_right_out;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__166_ccff_tail;
wire [0:63] cbx_1__0__166_chanx_left_out;
wire [0:63] cbx_1__0__166_chanx_right_out;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__167_ccff_tail;
wire [0:63] cbx_1__0__167_chanx_left_out;
wire [0:63] cbx_1__0__167_chanx_right_out;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__168_ccff_tail;
wire [0:63] cbx_1__0__168_chanx_left_out;
wire [0:63] cbx_1__0__168_chanx_right_out;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__169_ccff_tail;
wire [0:63] cbx_1__0__169_chanx_left_out;
wire [0:63] cbx_1__0__169_chanx_right_out;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__16_ccff_tail;
wire [0:63] cbx_1__0__16_chanx_left_out;
wire [0:63] cbx_1__0__16_chanx_right_out;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__170_ccff_tail;
wire [0:63] cbx_1__0__170_chanx_left_out;
wire [0:63] cbx_1__0__170_chanx_right_out;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__171_ccff_tail;
wire [0:63] cbx_1__0__171_chanx_left_out;
wire [0:63] cbx_1__0__171_chanx_right_out;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__172_ccff_tail;
wire [0:63] cbx_1__0__172_chanx_left_out;
wire [0:63] cbx_1__0__172_chanx_right_out;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__173_ccff_tail;
wire [0:63] cbx_1__0__173_chanx_left_out;
wire [0:63] cbx_1__0__173_chanx_right_out;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__174_ccff_tail;
wire [0:63] cbx_1__0__174_chanx_left_out;
wire [0:63] cbx_1__0__174_chanx_right_out;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__175_ccff_tail;
wire [0:63] cbx_1__0__175_chanx_left_out;
wire [0:63] cbx_1__0__175_chanx_right_out;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__176_ccff_tail;
wire [0:63] cbx_1__0__176_chanx_left_out;
wire [0:63] cbx_1__0__176_chanx_right_out;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__177_ccff_tail;
wire [0:63] cbx_1__0__177_chanx_left_out;
wire [0:63] cbx_1__0__177_chanx_right_out;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__178_ccff_tail;
wire [0:63] cbx_1__0__178_chanx_left_out;
wire [0:63] cbx_1__0__178_chanx_right_out;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__179_ccff_tail;
wire [0:63] cbx_1__0__179_chanx_left_out;
wire [0:63] cbx_1__0__179_chanx_right_out;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__17_ccff_tail;
wire [0:63] cbx_1__0__17_chanx_left_out;
wire [0:63] cbx_1__0__17_chanx_right_out;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__180_ccff_tail;
wire [0:63] cbx_1__0__180_chanx_left_out;
wire [0:63] cbx_1__0__180_chanx_right_out;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__181_ccff_tail;
wire [0:63] cbx_1__0__181_chanx_left_out;
wire [0:63] cbx_1__0__181_chanx_right_out;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__182_ccff_tail;
wire [0:63] cbx_1__0__182_chanx_left_out;
wire [0:63] cbx_1__0__182_chanx_right_out;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__183_ccff_tail;
wire [0:63] cbx_1__0__183_chanx_left_out;
wire [0:63] cbx_1__0__183_chanx_right_out;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__184_ccff_tail;
wire [0:63] cbx_1__0__184_chanx_left_out;
wire [0:63] cbx_1__0__184_chanx_right_out;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__185_ccff_tail;
wire [0:63] cbx_1__0__185_chanx_left_out;
wire [0:63] cbx_1__0__185_chanx_right_out;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__186_ccff_tail;
wire [0:63] cbx_1__0__186_chanx_left_out;
wire [0:63] cbx_1__0__186_chanx_right_out;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__187_ccff_tail;
wire [0:63] cbx_1__0__187_chanx_left_out;
wire [0:63] cbx_1__0__187_chanx_right_out;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__188_ccff_tail;
wire [0:63] cbx_1__0__188_chanx_left_out;
wire [0:63] cbx_1__0__188_chanx_right_out;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__189_ccff_tail;
wire [0:63] cbx_1__0__189_chanx_left_out;
wire [0:63] cbx_1__0__189_chanx_right_out;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__18_ccff_tail;
wire [0:63] cbx_1__0__18_chanx_left_out;
wire [0:63] cbx_1__0__18_chanx_right_out;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__190_ccff_tail;
wire [0:63] cbx_1__0__190_chanx_left_out;
wire [0:63] cbx_1__0__190_chanx_right_out;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__191_ccff_tail;
wire [0:63] cbx_1__0__191_chanx_left_out;
wire [0:63] cbx_1__0__191_chanx_right_out;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__192_ccff_tail;
wire [0:63] cbx_1__0__192_chanx_left_out;
wire [0:63] cbx_1__0__192_chanx_right_out;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__193_ccff_tail;
wire [0:63] cbx_1__0__193_chanx_left_out;
wire [0:63] cbx_1__0__193_chanx_right_out;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__194_ccff_tail;
wire [0:63] cbx_1__0__194_chanx_left_out;
wire [0:63] cbx_1__0__194_chanx_right_out;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__195_ccff_tail;
wire [0:63] cbx_1__0__195_chanx_left_out;
wire [0:63] cbx_1__0__195_chanx_right_out;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__196_ccff_tail;
wire [0:63] cbx_1__0__196_chanx_left_out;
wire [0:63] cbx_1__0__196_chanx_right_out;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__197_ccff_tail;
wire [0:63] cbx_1__0__197_chanx_left_out;
wire [0:63] cbx_1__0__197_chanx_right_out;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__198_ccff_tail;
wire [0:63] cbx_1__0__198_chanx_left_out;
wire [0:63] cbx_1__0__198_chanx_right_out;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__199_ccff_tail;
wire [0:63] cbx_1__0__199_chanx_left_out;
wire [0:63] cbx_1__0__199_chanx_right_out;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__19_ccff_tail;
wire [0:63] cbx_1__0__19_chanx_left_out;
wire [0:63] cbx_1__0__19_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:63] cbx_1__0__1_chanx_left_out;
wire [0:63] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__200_ccff_tail;
wire [0:63] cbx_1__0__200_chanx_left_out;
wire [0:63] cbx_1__0__200_chanx_right_out;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__201_ccff_tail;
wire [0:63] cbx_1__0__201_chanx_left_out;
wire [0:63] cbx_1__0__201_chanx_right_out;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__202_ccff_tail;
wire [0:63] cbx_1__0__202_chanx_left_out;
wire [0:63] cbx_1__0__202_chanx_right_out;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__203_ccff_tail;
wire [0:63] cbx_1__0__203_chanx_left_out;
wire [0:63] cbx_1__0__203_chanx_right_out;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__204_ccff_tail;
wire [0:63] cbx_1__0__204_chanx_left_out;
wire [0:63] cbx_1__0__204_chanx_right_out;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__205_ccff_tail;
wire [0:63] cbx_1__0__205_chanx_left_out;
wire [0:63] cbx_1__0__205_chanx_right_out;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__206_ccff_tail;
wire [0:63] cbx_1__0__206_chanx_left_out;
wire [0:63] cbx_1__0__206_chanx_right_out;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__207_ccff_tail;
wire [0:63] cbx_1__0__207_chanx_left_out;
wire [0:63] cbx_1__0__207_chanx_right_out;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__208_ccff_tail;
wire [0:63] cbx_1__0__208_chanx_left_out;
wire [0:63] cbx_1__0__208_chanx_right_out;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__209_ccff_tail;
wire [0:63] cbx_1__0__209_chanx_left_out;
wire [0:63] cbx_1__0__209_chanx_right_out;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__20_ccff_tail;
wire [0:63] cbx_1__0__20_chanx_left_out;
wire [0:63] cbx_1__0__20_chanx_right_out;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__210_ccff_tail;
wire [0:63] cbx_1__0__210_chanx_left_out;
wire [0:63] cbx_1__0__210_chanx_right_out;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__211_ccff_tail;
wire [0:63] cbx_1__0__211_chanx_left_out;
wire [0:63] cbx_1__0__211_chanx_right_out;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__212_ccff_tail;
wire [0:63] cbx_1__0__212_chanx_left_out;
wire [0:63] cbx_1__0__212_chanx_right_out;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__213_ccff_tail;
wire [0:63] cbx_1__0__213_chanx_left_out;
wire [0:63] cbx_1__0__213_chanx_right_out;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__214_ccff_tail;
wire [0:63] cbx_1__0__214_chanx_left_out;
wire [0:63] cbx_1__0__214_chanx_right_out;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__215_ccff_tail;
wire [0:63] cbx_1__0__215_chanx_left_out;
wire [0:63] cbx_1__0__215_chanx_right_out;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__21_ccff_tail;
wire [0:63] cbx_1__0__21_chanx_left_out;
wire [0:63] cbx_1__0__21_chanx_right_out;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__22_ccff_tail;
wire [0:63] cbx_1__0__22_chanx_left_out;
wire [0:63] cbx_1__0__22_chanx_right_out;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__23_ccff_tail;
wire [0:63] cbx_1__0__23_chanx_left_out;
wire [0:63] cbx_1__0__23_chanx_right_out;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__24_ccff_tail;
wire [0:63] cbx_1__0__24_chanx_left_out;
wire [0:63] cbx_1__0__24_chanx_right_out;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__25_ccff_tail;
wire [0:63] cbx_1__0__25_chanx_left_out;
wire [0:63] cbx_1__0__25_chanx_right_out;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__26_ccff_tail;
wire [0:63] cbx_1__0__26_chanx_left_out;
wire [0:63] cbx_1__0__26_chanx_right_out;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__27_ccff_tail;
wire [0:63] cbx_1__0__27_chanx_left_out;
wire [0:63] cbx_1__0__27_chanx_right_out;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__28_ccff_tail;
wire [0:63] cbx_1__0__28_chanx_left_out;
wire [0:63] cbx_1__0__28_chanx_right_out;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__29_ccff_tail;
wire [0:63] cbx_1__0__29_chanx_left_out;
wire [0:63] cbx_1__0__29_chanx_right_out;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:63] cbx_1__0__2_chanx_left_out;
wire [0:63] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__30_ccff_tail;
wire [0:63] cbx_1__0__30_chanx_left_out;
wire [0:63] cbx_1__0__30_chanx_right_out;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__31_ccff_tail;
wire [0:63] cbx_1__0__31_chanx_left_out;
wire [0:63] cbx_1__0__31_chanx_right_out;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__32_ccff_tail;
wire [0:63] cbx_1__0__32_chanx_left_out;
wire [0:63] cbx_1__0__32_chanx_right_out;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__33_ccff_tail;
wire [0:63] cbx_1__0__33_chanx_left_out;
wire [0:63] cbx_1__0__33_chanx_right_out;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__34_ccff_tail;
wire [0:63] cbx_1__0__34_chanx_left_out;
wire [0:63] cbx_1__0__34_chanx_right_out;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__35_ccff_tail;
wire [0:63] cbx_1__0__35_chanx_left_out;
wire [0:63] cbx_1__0__35_chanx_right_out;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__36_ccff_tail;
wire [0:63] cbx_1__0__36_chanx_left_out;
wire [0:63] cbx_1__0__36_chanx_right_out;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__37_ccff_tail;
wire [0:63] cbx_1__0__37_chanx_left_out;
wire [0:63] cbx_1__0__37_chanx_right_out;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__38_ccff_tail;
wire [0:63] cbx_1__0__38_chanx_left_out;
wire [0:63] cbx_1__0__38_chanx_right_out;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__39_ccff_tail;
wire [0:63] cbx_1__0__39_chanx_left_out;
wire [0:63] cbx_1__0__39_chanx_right_out;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:63] cbx_1__0__3_chanx_left_out;
wire [0:63] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__40_ccff_tail;
wire [0:63] cbx_1__0__40_chanx_left_out;
wire [0:63] cbx_1__0__40_chanx_right_out;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__41_ccff_tail;
wire [0:63] cbx_1__0__41_chanx_left_out;
wire [0:63] cbx_1__0__41_chanx_right_out;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__42_ccff_tail;
wire [0:63] cbx_1__0__42_chanx_left_out;
wire [0:63] cbx_1__0__42_chanx_right_out;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__43_ccff_tail;
wire [0:63] cbx_1__0__43_chanx_left_out;
wire [0:63] cbx_1__0__43_chanx_right_out;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__44_ccff_tail;
wire [0:63] cbx_1__0__44_chanx_left_out;
wire [0:63] cbx_1__0__44_chanx_right_out;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__45_ccff_tail;
wire [0:63] cbx_1__0__45_chanx_left_out;
wire [0:63] cbx_1__0__45_chanx_right_out;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__46_ccff_tail;
wire [0:63] cbx_1__0__46_chanx_left_out;
wire [0:63] cbx_1__0__46_chanx_right_out;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__47_ccff_tail;
wire [0:63] cbx_1__0__47_chanx_left_out;
wire [0:63] cbx_1__0__47_chanx_right_out;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__48_ccff_tail;
wire [0:63] cbx_1__0__48_chanx_left_out;
wire [0:63] cbx_1__0__48_chanx_right_out;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__49_ccff_tail;
wire [0:63] cbx_1__0__49_chanx_left_out;
wire [0:63] cbx_1__0__49_chanx_right_out;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:63] cbx_1__0__4_chanx_left_out;
wire [0:63] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__50_ccff_tail;
wire [0:63] cbx_1__0__50_chanx_left_out;
wire [0:63] cbx_1__0__50_chanx_right_out;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__51_ccff_tail;
wire [0:63] cbx_1__0__51_chanx_left_out;
wire [0:63] cbx_1__0__51_chanx_right_out;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__52_ccff_tail;
wire [0:63] cbx_1__0__52_chanx_left_out;
wire [0:63] cbx_1__0__52_chanx_right_out;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__53_ccff_tail;
wire [0:63] cbx_1__0__53_chanx_left_out;
wire [0:63] cbx_1__0__53_chanx_right_out;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__54_ccff_tail;
wire [0:63] cbx_1__0__54_chanx_left_out;
wire [0:63] cbx_1__0__54_chanx_right_out;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__55_ccff_tail;
wire [0:63] cbx_1__0__55_chanx_left_out;
wire [0:63] cbx_1__0__55_chanx_right_out;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__56_ccff_tail;
wire [0:63] cbx_1__0__56_chanx_left_out;
wire [0:63] cbx_1__0__56_chanx_right_out;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__57_ccff_tail;
wire [0:63] cbx_1__0__57_chanx_left_out;
wire [0:63] cbx_1__0__57_chanx_right_out;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__58_ccff_tail;
wire [0:63] cbx_1__0__58_chanx_left_out;
wire [0:63] cbx_1__0__58_chanx_right_out;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__59_ccff_tail;
wire [0:63] cbx_1__0__59_chanx_left_out;
wire [0:63] cbx_1__0__59_chanx_right_out;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:63] cbx_1__0__5_chanx_left_out;
wire [0:63] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__60_ccff_tail;
wire [0:63] cbx_1__0__60_chanx_left_out;
wire [0:63] cbx_1__0__60_chanx_right_out;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__61_ccff_tail;
wire [0:63] cbx_1__0__61_chanx_left_out;
wire [0:63] cbx_1__0__61_chanx_right_out;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__62_ccff_tail;
wire [0:63] cbx_1__0__62_chanx_left_out;
wire [0:63] cbx_1__0__62_chanx_right_out;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__63_ccff_tail;
wire [0:63] cbx_1__0__63_chanx_left_out;
wire [0:63] cbx_1__0__63_chanx_right_out;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__64_ccff_tail;
wire [0:63] cbx_1__0__64_chanx_left_out;
wire [0:63] cbx_1__0__64_chanx_right_out;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__65_ccff_tail;
wire [0:63] cbx_1__0__65_chanx_left_out;
wire [0:63] cbx_1__0__65_chanx_right_out;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__66_ccff_tail;
wire [0:63] cbx_1__0__66_chanx_left_out;
wire [0:63] cbx_1__0__66_chanx_right_out;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__67_ccff_tail;
wire [0:63] cbx_1__0__67_chanx_left_out;
wire [0:63] cbx_1__0__67_chanx_right_out;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__68_ccff_tail;
wire [0:63] cbx_1__0__68_chanx_left_out;
wire [0:63] cbx_1__0__68_chanx_right_out;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__69_ccff_tail;
wire [0:63] cbx_1__0__69_chanx_left_out;
wire [0:63] cbx_1__0__69_chanx_right_out;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:63] cbx_1__0__6_chanx_left_out;
wire [0:63] cbx_1__0__6_chanx_right_out;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__70_ccff_tail;
wire [0:63] cbx_1__0__70_chanx_left_out;
wire [0:63] cbx_1__0__70_chanx_right_out;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__71_ccff_tail;
wire [0:63] cbx_1__0__71_chanx_left_out;
wire [0:63] cbx_1__0__71_chanx_right_out;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__72_ccff_tail;
wire [0:63] cbx_1__0__72_chanx_left_out;
wire [0:63] cbx_1__0__72_chanx_right_out;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__73_ccff_tail;
wire [0:63] cbx_1__0__73_chanx_left_out;
wire [0:63] cbx_1__0__73_chanx_right_out;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__74_ccff_tail;
wire [0:63] cbx_1__0__74_chanx_left_out;
wire [0:63] cbx_1__0__74_chanx_right_out;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__75_ccff_tail;
wire [0:63] cbx_1__0__75_chanx_left_out;
wire [0:63] cbx_1__0__75_chanx_right_out;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__76_ccff_tail;
wire [0:63] cbx_1__0__76_chanx_left_out;
wire [0:63] cbx_1__0__76_chanx_right_out;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__77_ccff_tail;
wire [0:63] cbx_1__0__77_chanx_left_out;
wire [0:63] cbx_1__0__77_chanx_right_out;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__78_ccff_tail;
wire [0:63] cbx_1__0__78_chanx_left_out;
wire [0:63] cbx_1__0__78_chanx_right_out;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__79_ccff_tail;
wire [0:63] cbx_1__0__79_chanx_left_out;
wire [0:63] cbx_1__0__79_chanx_right_out;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__7_ccff_tail;
wire [0:63] cbx_1__0__7_chanx_left_out;
wire [0:63] cbx_1__0__7_chanx_right_out;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__80_ccff_tail;
wire [0:63] cbx_1__0__80_chanx_left_out;
wire [0:63] cbx_1__0__80_chanx_right_out;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__81_ccff_tail;
wire [0:63] cbx_1__0__81_chanx_left_out;
wire [0:63] cbx_1__0__81_chanx_right_out;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__82_ccff_tail;
wire [0:63] cbx_1__0__82_chanx_left_out;
wire [0:63] cbx_1__0__82_chanx_right_out;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__83_ccff_tail;
wire [0:63] cbx_1__0__83_chanx_left_out;
wire [0:63] cbx_1__0__83_chanx_right_out;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__84_ccff_tail;
wire [0:63] cbx_1__0__84_chanx_left_out;
wire [0:63] cbx_1__0__84_chanx_right_out;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__85_ccff_tail;
wire [0:63] cbx_1__0__85_chanx_left_out;
wire [0:63] cbx_1__0__85_chanx_right_out;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__86_ccff_tail;
wire [0:63] cbx_1__0__86_chanx_left_out;
wire [0:63] cbx_1__0__86_chanx_right_out;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__87_ccff_tail;
wire [0:63] cbx_1__0__87_chanx_left_out;
wire [0:63] cbx_1__0__87_chanx_right_out;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__88_ccff_tail;
wire [0:63] cbx_1__0__88_chanx_left_out;
wire [0:63] cbx_1__0__88_chanx_right_out;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__89_ccff_tail;
wire [0:63] cbx_1__0__89_chanx_left_out;
wire [0:63] cbx_1__0__89_chanx_right_out;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__8_ccff_tail;
wire [0:63] cbx_1__0__8_chanx_left_out;
wire [0:63] cbx_1__0__8_chanx_right_out;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__90_ccff_tail;
wire [0:63] cbx_1__0__90_chanx_left_out;
wire [0:63] cbx_1__0__90_chanx_right_out;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__91_ccff_tail;
wire [0:63] cbx_1__0__91_chanx_left_out;
wire [0:63] cbx_1__0__91_chanx_right_out;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__92_ccff_tail;
wire [0:63] cbx_1__0__92_chanx_left_out;
wire [0:63] cbx_1__0__92_chanx_right_out;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__93_ccff_tail;
wire [0:63] cbx_1__0__93_chanx_left_out;
wire [0:63] cbx_1__0__93_chanx_right_out;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__94_ccff_tail;
wire [0:63] cbx_1__0__94_chanx_left_out;
wire [0:63] cbx_1__0__94_chanx_right_out;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__95_ccff_tail;
wire [0:63] cbx_1__0__95_chanx_left_out;
wire [0:63] cbx_1__0__95_chanx_right_out;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__96_ccff_tail;
wire [0:63] cbx_1__0__96_chanx_left_out;
wire [0:63] cbx_1__0__96_chanx_right_out;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__97_ccff_tail;
wire [0:63] cbx_1__0__97_chanx_left_out;
wire [0:63] cbx_1__0__97_chanx_right_out;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__98_ccff_tail;
wire [0:63] cbx_1__0__98_chanx_left_out;
wire [0:63] cbx_1__0__98_chanx_right_out;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__99_ccff_tail;
wire [0:63] cbx_1__0__99_chanx_left_out;
wire [0:63] cbx_1__0__99_chanx_right_out;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__9_ccff_tail;
wire [0:63] cbx_1__0__9_chanx_left_out;
wire [0:63] cbx_1__0__9_chanx_right_out;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__0_ccff_tail;
wire [0:63] cbx_1__18__0_chanx_left_out;
wire [0:63] cbx_1__18__0_chanx_right_out;
wire [0:0] cbx_1__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__10_ccff_tail;
wire [0:63] cbx_1__18__10_chanx_left_out;
wire [0:63] cbx_1__18__10_chanx_right_out;
wire [0:0] cbx_1__18__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__11_ccff_tail;
wire [0:63] cbx_1__18__11_chanx_left_out;
wire [0:63] cbx_1__18__11_chanx_right_out;
wire [0:0] cbx_1__18__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__1_ccff_tail;
wire [0:63] cbx_1__18__1_chanx_left_out;
wire [0:63] cbx_1__18__1_chanx_right_out;
wire [0:0] cbx_1__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__2_ccff_tail;
wire [0:63] cbx_1__18__2_chanx_left_out;
wire [0:63] cbx_1__18__2_chanx_right_out;
wire [0:0] cbx_1__18__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__3_ccff_tail;
wire [0:63] cbx_1__18__3_chanx_left_out;
wire [0:63] cbx_1__18__3_chanx_right_out;
wire [0:0] cbx_1__18__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__4_ccff_tail;
wire [0:63] cbx_1__18__4_chanx_left_out;
wire [0:63] cbx_1__18__4_chanx_right_out;
wire [0:0] cbx_1__18__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__5_ccff_tail;
wire [0:63] cbx_1__18__5_chanx_left_out;
wire [0:63] cbx_1__18__5_chanx_right_out;
wire [0:0] cbx_1__18__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__6_ccff_tail;
wire [0:63] cbx_1__18__6_chanx_left_out;
wire [0:63] cbx_1__18__6_chanx_right_out;
wire [0:0] cbx_1__18__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__7_ccff_tail;
wire [0:63] cbx_1__18__7_chanx_left_out;
wire [0:63] cbx_1__18__7_chanx_right_out;
wire [0:0] cbx_1__18__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__8_ccff_tail;
wire [0:63] cbx_1__18__8_chanx_left_out;
wire [0:63] cbx_1__18__8_chanx_right_out;
wire [0:0] cbx_1__18__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__18__9_ccff_tail;
wire [0:63] cbx_1__18__9_chanx_left_out;
wire [0:63] cbx_1__18__9_chanx_right_out;
wire [0:0] cbx_1__18__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_4__0__0_ccff_tail;
wire [0:63] cbx_4__0__0_chanx_left_out;
wire [0:63] cbx_4__0__0_chanx_right_out;
wire [0:0] cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_4__0__1_ccff_tail;
wire [0:63] cbx_4__0__1_chanx_left_out;
wire [0:63] cbx_4__0__1_chanx_right_out;
wire [0:0] cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__18__0_ccff_tail;
wire [0:63] cbx_4__18__0_chanx_left_out;
wire [0:63] cbx_4__18__0_chanx_right_out;
wire [0:0] cbx_4__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__18__1_ccff_tail;
wire [0:63] cbx_4__18__1_chanx_left_out;
wire [0:63] cbx_4__18__1_chanx_right_out;
wire [0:0] cbx_4__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__0_ccff_tail;
wire [0:63] cbx_4__1__0_chanx_left_out;
wire [0:63] cbx_4__1__0_chanx_right_out;
wire [0:0] cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__10_ccff_tail;
wire [0:63] cbx_4__1__10_chanx_left_out;
wire [0:63] cbx_4__1__10_chanx_right_out;
wire [0:0] cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__11_ccff_tail;
wire [0:63] cbx_4__1__11_chanx_left_out;
wire [0:63] cbx_4__1__11_chanx_right_out;
wire [0:0] cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__12_ccff_tail;
wire [0:63] cbx_4__1__12_chanx_left_out;
wire [0:63] cbx_4__1__12_chanx_right_out;
wire [0:0] cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__13_ccff_tail;
wire [0:63] cbx_4__1__13_chanx_left_out;
wire [0:63] cbx_4__1__13_chanx_right_out;
wire [0:0] cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__14_ccff_tail;
wire [0:63] cbx_4__1__14_chanx_left_out;
wire [0:63] cbx_4__1__14_chanx_right_out;
wire [0:0] cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__15_ccff_tail;
wire [0:63] cbx_4__1__15_chanx_left_out;
wire [0:63] cbx_4__1__15_chanx_right_out;
wire [0:0] cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__16_ccff_tail;
wire [0:63] cbx_4__1__16_chanx_left_out;
wire [0:63] cbx_4__1__16_chanx_right_out;
wire [0:0] cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__17_ccff_tail;
wire [0:63] cbx_4__1__17_chanx_left_out;
wire [0:63] cbx_4__1__17_chanx_right_out;
wire [0:0] cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__1_ccff_tail;
wire [0:63] cbx_4__1__1_chanx_left_out;
wire [0:63] cbx_4__1__1_chanx_right_out;
wire [0:0] cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__2_ccff_tail;
wire [0:63] cbx_4__1__2_chanx_left_out;
wire [0:63] cbx_4__1__2_chanx_right_out;
wire [0:0] cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__3_ccff_tail;
wire [0:63] cbx_4__1__3_chanx_left_out;
wire [0:63] cbx_4__1__3_chanx_right_out;
wire [0:0] cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__4_ccff_tail;
wire [0:63] cbx_4__1__4_chanx_left_out;
wire [0:63] cbx_4__1__4_chanx_right_out;
wire [0:0] cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__5_ccff_tail;
wire [0:63] cbx_4__1__5_chanx_left_out;
wire [0:63] cbx_4__1__5_chanx_right_out;
wire [0:0] cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__6_ccff_tail;
wire [0:63] cbx_4__1__6_chanx_left_out;
wire [0:63] cbx_4__1__6_chanx_right_out;
wire [0:0] cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__7_ccff_tail;
wire [0:63] cbx_4__1__7_chanx_left_out;
wire [0:63] cbx_4__1__7_chanx_right_out;
wire [0:0] cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__8_ccff_tail;
wire [0:63] cbx_4__1__8_chanx_left_out;
wire [0:63] cbx_4__1__8_chanx_right_out;
wire [0:0] cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_4__1__9_ccff_tail;
wire [0:63] cbx_4__1__9_chanx_left_out;
wire [0:63] cbx_4__1__9_chanx_right_out;
wire [0:0] cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_;
wire [0:0] cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_;
wire [0:0] cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_;
wire [0:0] cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__0_ccff_tail;
wire [0:63] cbx_4__2__0_chanx_left_out;
wire [0:63] cbx_4__2__0_chanx_right_out;
wire [0:0] cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__10_ccff_tail;
wire [0:63] cbx_4__2__10_chanx_left_out;
wire [0:63] cbx_4__2__10_chanx_right_out;
wire [0:0] cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__11_ccff_tail;
wire [0:63] cbx_4__2__11_chanx_left_out;
wire [0:63] cbx_4__2__11_chanx_right_out;
wire [0:0] cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__12_ccff_tail;
wire [0:63] cbx_4__2__12_chanx_left_out;
wire [0:63] cbx_4__2__12_chanx_right_out;
wire [0:0] cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__13_ccff_tail;
wire [0:63] cbx_4__2__13_chanx_left_out;
wire [0:63] cbx_4__2__13_chanx_right_out;
wire [0:0] cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__14_ccff_tail;
wire [0:63] cbx_4__2__14_chanx_left_out;
wire [0:63] cbx_4__2__14_chanx_right_out;
wire [0:0] cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__15_ccff_tail;
wire [0:63] cbx_4__2__15_chanx_left_out;
wire [0:63] cbx_4__2__15_chanx_right_out;
wire [0:0] cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__1_ccff_tail;
wire [0:63] cbx_4__2__1_chanx_left_out;
wire [0:63] cbx_4__2__1_chanx_right_out;
wire [0:0] cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__2_ccff_tail;
wire [0:63] cbx_4__2__2_chanx_left_out;
wire [0:63] cbx_4__2__2_chanx_right_out;
wire [0:0] cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__3_ccff_tail;
wire [0:63] cbx_4__2__3_chanx_left_out;
wire [0:63] cbx_4__2__3_chanx_right_out;
wire [0:0] cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__4_ccff_tail;
wire [0:63] cbx_4__2__4_chanx_left_out;
wire [0:63] cbx_4__2__4_chanx_right_out;
wire [0:0] cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__5_ccff_tail;
wire [0:63] cbx_4__2__5_chanx_left_out;
wire [0:63] cbx_4__2__5_chanx_right_out;
wire [0:0] cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__6_ccff_tail;
wire [0:63] cbx_4__2__6_chanx_left_out;
wire [0:63] cbx_4__2__6_chanx_right_out;
wire [0:0] cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__7_ccff_tail;
wire [0:63] cbx_4__2__7_chanx_left_out;
wire [0:63] cbx_4__2__7_chanx_right_out;
wire [0:0] cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__8_ccff_tail;
wire [0:63] cbx_4__2__8_chanx_left_out;
wire [0:63] cbx_4__2__8_chanx_right_out;
wire [0:0] cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_;
wire [0:0] cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_;
wire [0:0] cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_;
wire [0:0] cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_;
wire [0:0] cbx_4__2__9_ccff_tail;
wire [0:63] cbx_4__2__9_chanx_left_out;
wire [0:63] cbx_4__2__9_chanx_right_out;
wire [0:0] cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:63] cby_0__1__0_chany_bottom_out;
wire [0:63] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__10_ccff_tail;
wire [0:63] cby_0__1__10_chany_bottom_out;
wire [0:63] cby_0__1__10_chany_top_out;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__11_ccff_tail;
wire [0:63] cby_0__1__11_chany_bottom_out;
wire [0:63] cby_0__1__11_chany_top_out;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__12_ccff_tail;
wire [0:63] cby_0__1__12_chany_bottom_out;
wire [0:63] cby_0__1__12_chany_top_out;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__13_ccff_tail;
wire [0:63] cby_0__1__13_chany_bottom_out;
wire [0:63] cby_0__1__13_chany_top_out;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__14_ccff_tail;
wire [0:63] cby_0__1__14_chany_bottom_out;
wire [0:63] cby_0__1__14_chany_top_out;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__15_ccff_tail;
wire [0:63] cby_0__1__15_chany_bottom_out;
wire [0:63] cby_0__1__15_chany_top_out;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__16_ccff_tail;
wire [0:63] cby_0__1__16_chany_bottom_out;
wire [0:63] cby_0__1__16_chany_top_out;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__17_ccff_tail;
wire [0:63] cby_0__1__17_chany_bottom_out;
wire [0:63] cby_0__1__17_chany_top_out;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:63] cby_0__1__1_chany_bottom_out;
wire [0:63] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:63] cby_0__1__2_chany_bottom_out;
wire [0:63] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:63] cby_0__1__3_chany_bottom_out;
wire [0:63] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:63] cby_0__1__4_chany_bottom_out;
wire [0:63] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__5_ccff_tail;
wire [0:63] cby_0__1__5_chany_bottom_out;
wire [0:63] cby_0__1__5_chany_top_out;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__6_ccff_tail;
wire [0:63] cby_0__1__6_chany_bottom_out;
wire [0:63] cby_0__1__6_chany_top_out;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__7_ccff_tail;
wire [0:63] cby_0__1__7_chany_bottom_out;
wire [0:63] cby_0__1__7_chany_top_out;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__8_ccff_tail;
wire [0:63] cby_0__1__8_chany_bottom_out;
wire [0:63] cby_0__1__8_chany_top_out;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__9_ccff_tail;
wire [0:63] cby_0__1__9_chany_bottom_out;
wire [0:63] cby_0__1__9_chany_top_out;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:63] cby_14__1__0_chany_bottom_out;
wire [0:63] cby_14__1__0_chany_top_out;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__10_ccff_tail;
wire [0:63] cby_14__1__10_chany_bottom_out;
wire [0:63] cby_14__1__10_chany_top_out;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__11_ccff_tail;
wire [0:63] cby_14__1__11_chany_bottom_out;
wire [0:63] cby_14__1__11_chany_top_out;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__12_ccff_tail;
wire [0:63] cby_14__1__12_chany_bottom_out;
wire [0:63] cby_14__1__12_chany_top_out;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__13_ccff_tail;
wire [0:63] cby_14__1__13_chany_bottom_out;
wire [0:63] cby_14__1__13_chany_top_out;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__14_ccff_tail;
wire [0:63] cby_14__1__14_chany_bottom_out;
wire [0:63] cby_14__1__14_chany_top_out;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__15_ccff_tail;
wire [0:63] cby_14__1__15_chany_bottom_out;
wire [0:63] cby_14__1__15_chany_top_out;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__16_ccff_tail;
wire [0:63] cby_14__1__16_chany_bottom_out;
wire [0:63] cby_14__1__16_chany_top_out;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__17_ccff_tail;
wire [0:63] cby_14__1__17_chany_bottom_out;
wire [0:63] cby_14__1__17_chany_top_out;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__1_ccff_tail;
wire [0:63] cby_14__1__1_chany_bottom_out;
wire [0:63] cby_14__1__1_chany_top_out;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__2_ccff_tail;
wire [0:63] cby_14__1__2_chany_bottom_out;
wire [0:63] cby_14__1__2_chany_top_out;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__3_ccff_tail;
wire [0:63] cby_14__1__3_chany_bottom_out;
wire [0:63] cby_14__1__3_chany_top_out;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__4_ccff_tail;
wire [0:63] cby_14__1__4_chany_bottom_out;
wire [0:63] cby_14__1__4_chany_top_out;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__5_ccff_tail;
wire [0:63] cby_14__1__5_chany_bottom_out;
wire [0:63] cby_14__1__5_chany_top_out;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__6_ccff_tail;
wire [0:63] cby_14__1__6_chany_bottom_out;
wire [0:63] cby_14__1__6_chany_top_out;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__7_ccff_tail;
wire [0:63] cby_14__1__7_chany_bottom_out;
wire [0:63] cby_14__1__7_chany_top_out;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__8_ccff_tail;
wire [0:63] cby_14__1__8_chany_bottom_out;
wire [0:63] cby_14__1__8_chany_top_out;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_14__1__9_ccff_tail;
wire [0:63] cby_14__1__9_chany_bottom_out;
wire [0:63] cby_14__1__9_chany_top_out;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_14__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:63] cby_1__1__0_chany_bottom_out;
wire [0:63] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__100_ccff_tail;
wire [0:63] cby_1__1__100_chany_bottom_out;
wire [0:63] cby_1__1__100_chany_top_out;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__101_ccff_tail;
wire [0:63] cby_1__1__101_chany_bottom_out;
wire [0:63] cby_1__1__101_chany_top_out;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__102_ccff_tail;
wire [0:63] cby_1__1__102_chany_bottom_out;
wire [0:63] cby_1__1__102_chany_top_out;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__103_ccff_tail;
wire [0:63] cby_1__1__103_chany_bottom_out;
wire [0:63] cby_1__1__103_chany_top_out;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__104_ccff_tail;
wire [0:63] cby_1__1__104_chany_bottom_out;
wire [0:63] cby_1__1__104_chany_top_out;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__105_ccff_tail;
wire [0:63] cby_1__1__105_chany_bottom_out;
wire [0:63] cby_1__1__105_chany_top_out;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__106_ccff_tail;
wire [0:63] cby_1__1__106_chany_bottom_out;
wire [0:63] cby_1__1__106_chany_top_out;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__107_ccff_tail;
wire [0:63] cby_1__1__107_chany_bottom_out;
wire [0:63] cby_1__1__107_chany_top_out;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__108_ccff_tail;
wire [0:63] cby_1__1__108_chany_bottom_out;
wire [0:63] cby_1__1__108_chany_top_out;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__109_ccff_tail;
wire [0:63] cby_1__1__109_chany_bottom_out;
wire [0:63] cby_1__1__109_chany_top_out;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__10_ccff_tail;
wire [0:63] cby_1__1__10_chany_bottom_out;
wire [0:63] cby_1__1__10_chany_top_out;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__110_ccff_tail;
wire [0:63] cby_1__1__110_chany_bottom_out;
wire [0:63] cby_1__1__110_chany_top_out;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__111_ccff_tail;
wire [0:63] cby_1__1__111_chany_bottom_out;
wire [0:63] cby_1__1__111_chany_top_out;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__112_ccff_tail;
wire [0:63] cby_1__1__112_chany_bottom_out;
wire [0:63] cby_1__1__112_chany_top_out;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__113_ccff_tail;
wire [0:63] cby_1__1__113_chany_bottom_out;
wire [0:63] cby_1__1__113_chany_top_out;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__114_ccff_tail;
wire [0:63] cby_1__1__114_chany_bottom_out;
wire [0:63] cby_1__1__114_chany_top_out;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__115_ccff_tail;
wire [0:63] cby_1__1__115_chany_bottom_out;
wire [0:63] cby_1__1__115_chany_top_out;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__116_ccff_tail;
wire [0:63] cby_1__1__116_chany_bottom_out;
wire [0:63] cby_1__1__116_chany_top_out;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:63] cby_1__1__117_chany_bottom_out;
wire [0:63] cby_1__1__117_chany_top_out;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__118_ccff_tail;
wire [0:63] cby_1__1__118_chany_bottom_out;
wire [0:63] cby_1__1__118_chany_top_out;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__119_ccff_tail;
wire [0:63] cby_1__1__119_chany_bottom_out;
wire [0:63] cby_1__1__119_chany_top_out;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__11_ccff_tail;
wire [0:63] cby_1__1__11_chany_bottom_out;
wire [0:63] cby_1__1__11_chany_top_out;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__120_ccff_tail;
wire [0:63] cby_1__1__120_chany_bottom_out;
wire [0:63] cby_1__1__120_chany_top_out;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__121_ccff_tail;
wire [0:63] cby_1__1__121_chany_bottom_out;
wire [0:63] cby_1__1__121_chany_top_out;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__122_ccff_tail;
wire [0:63] cby_1__1__122_chany_bottom_out;
wire [0:63] cby_1__1__122_chany_top_out;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__123_ccff_tail;
wire [0:63] cby_1__1__123_chany_bottom_out;
wire [0:63] cby_1__1__123_chany_top_out;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__124_ccff_tail;
wire [0:63] cby_1__1__124_chany_bottom_out;
wire [0:63] cby_1__1__124_chany_top_out;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__125_ccff_tail;
wire [0:63] cby_1__1__125_chany_bottom_out;
wire [0:63] cby_1__1__125_chany_top_out;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__126_ccff_tail;
wire [0:63] cby_1__1__126_chany_bottom_out;
wire [0:63] cby_1__1__126_chany_top_out;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__127_ccff_tail;
wire [0:63] cby_1__1__127_chany_bottom_out;
wire [0:63] cby_1__1__127_chany_top_out;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__128_ccff_tail;
wire [0:63] cby_1__1__128_chany_bottom_out;
wire [0:63] cby_1__1__128_chany_top_out;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__129_ccff_tail;
wire [0:63] cby_1__1__129_chany_bottom_out;
wire [0:63] cby_1__1__129_chany_top_out;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__12_ccff_tail;
wire [0:63] cby_1__1__12_chany_bottom_out;
wire [0:63] cby_1__1__12_chany_top_out;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__130_ccff_tail;
wire [0:63] cby_1__1__130_chany_bottom_out;
wire [0:63] cby_1__1__130_chany_top_out;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__131_ccff_tail;
wire [0:63] cby_1__1__131_chany_bottom_out;
wire [0:63] cby_1__1__131_chany_top_out;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__132_ccff_tail;
wire [0:63] cby_1__1__132_chany_bottom_out;
wire [0:63] cby_1__1__132_chany_top_out;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__133_ccff_tail;
wire [0:63] cby_1__1__133_chany_bottom_out;
wire [0:63] cby_1__1__133_chany_top_out;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__134_ccff_tail;
wire [0:63] cby_1__1__134_chany_bottom_out;
wire [0:63] cby_1__1__134_chany_top_out;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__135_ccff_tail;
wire [0:63] cby_1__1__135_chany_bottom_out;
wire [0:63] cby_1__1__135_chany_top_out;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__136_ccff_tail;
wire [0:63] cby_1__1__136_chany_bottom_out;
wire [0:63] cby_1__1__136_chany_top_out;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__137_ccff_tail;
wire [0:63] cby_1__1__137_chany_bottom_out;
wire [0:63] cby_1__1__137_chany_top_out;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__138_ccff_tail;
wire [0:63] cby_1__1__138_chany_bottom_out;
wire [0:63] cby_1__1__138_chany_top_out;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__139_ccff_tail;
wire [0:63] cby_1__1__139_chany_bottom_out;
wire [0:63] cby_1__1__139_chany_top_out;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__13_ccff_tail;
wire [0:63] cby_1__1__13_chany_bottom_out;
wire [0:63] cby_1__1__13_chany_top_out;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__140_ccff_tail;
wire [0:63] cby_1__1__140_chany_bottom_out;
wire [0:63] cby_1__1__140_chany_top_out;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__141_ccff_tail;
wire [0:63] cby_1__1__141_chany_bottom_out;
wire [0:63] cby_1__1__141_chany_top_out;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__142_ccff_tail;
wire [0:63] cby_1__1__142_chany_bottom_out;
wire [0:63] cby_1__1__142_chany_top_out;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__143_ccff_tail;
wire [0:63] cby_1__1__143_chany_bottom_out;
wire [0:63] cby_1__1__143_chany_top_out;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__144_ccff_tail;
wire [0:63] cby_1__1__144_chany_bottom_out;
wire [0:63] cby_1__1__144_chany_top_out;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__145_ccff_tail;
wire [0:63] cby_1__1__145_chany_bottom_out;
wire [0:63] cby_1__1__145_chany_top_out;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__146_ccff_tail;
wire [0:63] cby_1__1__146_chany_bottom_out;
wire [0:63] cby_1__1__146_chany_top_out;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__147_ccff_tail;
wire [0:63] cby_1__1__147_chany_bottom_out;
wire [0:63] cby_1__1__147_chany_top_out;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__148_ccff_tail;
wire [0:63] cby_1__1__148_chany_bottom_out;
wire [0:63] cby_1__1__148_chany_top_out;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__149_ccff_tail;
wire [0:63] cby_1__1__149_chany_bottom_out;
wire [0:63] cby_1__1__149_chany_top_out;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__14_ccff_tail;
wire [0:63] cby_1__1__14_chany_bottom_out;
wire [0:63] cby_1__1__14_chany_top_out;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__150_ccff_tail;
wire [0:63] cby_1__1__150_chany_bottom_out;
wire [0:63] cby_1__1__150_chany_top_out;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__151_ccff_tail;
wire [0:63] cby_1__1__151_chany_bottom_out;
wire [0:63] cby_1__1__151_chany_top_out;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__152_ccff_tail;
wire [0:63] cby_1__1__152_chany_bottom_out;
wire [0:63] cby_1__1__152_chany_top_out;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__153_ccff_tail;
wire [0:63] cby_1__1__153_chany_bottom_out;
wire [0:63] cby_1__1__153_chany_top_out;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__154_ccff_tail;
wire [0:63] cby_1__1__154_chany_bottom_out;
wire [0:63] cby_1__1__154_chany_top_out;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__155_ccff_tail;
wire [0:63] cby_1__1__155_chany_bottom_out;
wire [0:63] cby_1__1__155_chany_top_out;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__156_ccff_tail;
wire [0:63] cby_1__1__156_chany_bottom_out;
wire [0:63] cby_1__1__156_chany_top_out;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__157_ccff_tail;
wire [0:63] cby_1__1__157_chany_bottom_out;
wire [0:63] cby_1__1__157_chany_top_out;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__158_ccff_tail;
wire [0:63] cby_1__1__158_chany_bottom_out;
wire [0:63] cby_1__1__158_chany_top_out;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__159_ccff_tail;
wire [0:63] cby_1__1__159_chany_bottom_out;
wire [0:63] cby_1__1__159_chany_top_out;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__15_ccff_tail;
wire [0:63] cby_1__1__15_chany_bottom_out;
wire [0:63] cby_1__1__15_chany_top_out;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__160_ccff_tail;
wire [0:63] cby_1__1__160_chany_bottom_out;
wire [0:63] cby_1__1__160_chany_top_out;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__161_ccff_tail;
wire [0:63] cby_1__1__161_chany_bottom_out;
wire [0:63] cby_1__1__161_chany_top_out;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__16_ccff_tail;
wire [0:63] cby_1__1__16_chany_bottom_out;
wire [0:63] cby_1__1__16_chany_top_out;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__17_ccff_tail;
wire [0:63] cby_1__1__17_chany_bottom_out;
wire [0:63] cby_1__1__17_chany_top_out;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__18_ccff_tail;
wire [0:63] cby_1__1__18_chany_bottom_out;
wire [0:63] cby_1__1__18_chany_top_out;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__19_ccff_tail;
wire [0:63] cby_1__1__19_chany_bottom_out;
wire [0:63] cby_1__1__19_chany_top_out;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:63] cby_1__1__1_chany_bottom_out;
wire [0:63] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__20_ccff_tail;
wire [0:63] cby_1__1__20_chany_bottom_out;
wire [0:63] cby_1__1__20_chany_top_out;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__21_ccff_tail;
wire [0:63] cby_1__1__21_chany_bottom_out;
wire [0:63] cby_1__1__21_chany_top_out;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__22_ccff_tail;
wire [0:63] cby_1__1__22_chany_bottom_out;
wire [0:63] cby_1__1__22_chany_top_out;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__23_ccff_tail;
wire [0:63] cby_1__1__23_chany_bottom_out;
wire [0:63] cby_1__1__23_chany_top_out;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__24_ccff_tail;
wire [0:63] cby_1__1__24_chany_bottom_out;
wire [0:63] cby_1__1__24_chany_top_out;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__25_ccff_tail;
wire [0:63] cby_1__1__25_chany_bottom_out;
wire [0:63] cby_1__1__25_chany_top_out;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__26_ccff_tail;
wire [0:63] cby_1__1__26_chany_bottom_out;
wire [0:63] cby_1__1__26_chany_top_out;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__27_ccff_tail;
wire [0:63] cby_1__1__27_chany_bottom_out;
wire [0:63] cby_1__1__27_chany_top_out;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__28_ccff_tail;
wire [0:63] cby_1__1__28_chany_bottom_out;
wire [0:63] cby_1__1__28_chany_top_out;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__29_ccff_tail;
wire [0:63] cby_1__1__29_chany_bottom_out;
wire [0:63] cby_1__1__29_chany_top_out;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__2_ccff_tail;
wire [0:63] cby_1__1__2_chany_bottom_out;
wire [0:63] cby_1__1__2_chany_top_out;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__30_ccff_tail;
wire [0:63] cby_1__1__30_chany_bottom_out;
wire [0:63] cby_1__1__30_chany_top_out;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__31_ccff_tail;
wire [0:63] cby_1__1__31_chany_bottom_out;
wire [0:63] cby_1__1__31_chany_top_out;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__32_ccff_tail;
wire [0:63] cby_1__1__32_chany_bottom_out;
wire [0:63] cby_1__1__32_chany_top_out;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__33_ccff_tail;
wire [0:63] cby_1__1__33_chany_bottom_out;
wire [0:63] cby_1__1__33_chany_top_out;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__34_ccff_tail;
wire [0:63] cby_1__1__34_chany_bottom_out;
wire [0:63] cby_1__1__34_chany_top_out;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__35_ccff_tail;
wire [0:63] cby_1__1__35_chany_bottom_out;
wire [0:63] cby_1__1__35_chany_top_out;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__36_ccff_tail;
wire [0:63] cby_1__1__36_chany_bottom_out;
wire [0:63] cby_1__1__36_chany_top_out;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__37_ccff_tail;
wire [0:63] cby_1__1__37_chany_bottom_out;
wire [0:63] cby_1__1__37_chany_top_out;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__38_ccff_tail;
wire [0:63] cby_1__1__38_chany_bottom_out;
wire [0:63] cby_1__1__38_chany_top_out;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__39_ccff_tail;
wire [0:63] cby_1__1__39_chany_bottom_out;
wire [0:63] cby_1__1__39_chany_top_out;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__3_ccff_tail;
wire [0:63] cby_1__1__3_chany_bottom_out;
wire [0:63] cby_1__1__3_chany_top_out;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__40_ccff_tail;
wire [0:63] cby_1__1__40_chany_bottom_out;
wire [0:63] cby_1__1__40_chany_top_out;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__41_ccff_tail;
wire [0:63] cby_1__1__41_chany_bottom_out;
wire [0:63] cby_1__1__41_chany_top_out;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__42_ccff_tail;
wire [0:63] cby_1__1__42_chany_bottom_out;
wire [0:63] cby_1__1__42_chany_top_out;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__43_ccff_tail;
wire [0:63] cby_1__1__43_chany_bottom_out;
wire [0:63] cby_1__1__43_chany_top_out;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__44_ccff_tail;
wire [0:63] cby_1__1__44_chany_bottom_out;
wire [0:63] cby_1__1__44_chany_top_out;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__45_ccff_tail;
wire [0:63] cby_1__1__45_chany_bottom_out;
wire [0:63] cby_1__1__45_chany_top_out;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__46_ccff_tail;
wire [0:63] cby_1__1__46_chany_bottom_out;
wire [0:63] cby_1__1__46_chany_top_out;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__47_ccff_tail;
wire [0:63] cby_1__1__47_chany_bottom_out;
wire [0:63] cby_1__1__47_chany_top_out;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__48_ccff_tail;
wire [0:63] cby_1__1__48_chany_bottom_out;
wire [0:63] cby_1__1__48_chany_top_out;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__49_ccff_tail;
wire [0:63] cby_1__1__49_chany_bottom_out;
wire [0:63] cby_1__1__49_chany_top_out;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__4_ccff_tail;
wire [0:63] cby_1__1__4_chany_bottom_out;
wire [0:63] cby_1__1__4_chany_top_out;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__50_ccff_tail;
wire [0:63] cby_1__1__50_chany_bottom_out;
wire [0:63] cby_1__1__50_chany_top_out;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__51_ccff_tail;
wire [0:63] cby_1__1__51_chany_bottom_out;
wire [0:63] cby_1__1__51_chany_top_out;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__52_ccff_tail;
wire [0:63] cby_1__1__52_chany_bottom_out;
wire [0:63] cby_1__1__52_chany_top_out;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__53_ccff_tail;
wire [0:63] cby_1__1__53_chany_bottom_out;
wire [0:63] cby_1__1__53_chany_top_out;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__54_ccff_tail;
wire [0:63] cby_1__1__54_chany_bottom_out;
wire [0:63] cby_1__1__54_chany_top_out;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__55_ccff_tail;
wire [0:63] cby_1__1__55_chany_bottom_out;
wire [0:63] cby_1__1__55_chany_top_out;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__56_ccff_tail;
wire [0:63] cby_1__1__56_chany_bottom_out;
wire [0:63] cby_1__1__56_chany_top_out;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__57_ccff_tail;
wire [0:63] cby_1__1__57_chany_bottom_out;
wire [0:63] cby_1__1__57_chany_top_out;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__58_ccff_tail;
wire [0:63] cby_1__1__58_chany_bottom_out;
wire [0:63] cby_1__1__58_chany_top_out;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__59_ccff_tail;
wire [0:63] cby_1__1__59_chany_bottom_out;
wire [0:63] cby_1__1__59_chany_top_out;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__5_ccff_tail;
wire [0:63] cby_1__1__5_chany_bottom_out;
wire [0:63] cby_1__1__5_chany_top_out;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__60_ccff_tail;
wire [0:63] cby_1__1__60_chany_bottom_out;
wire [0:63] cby_1__1__60_chany_top_out;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__61_ccff_tail;
wire [0:63] cby_1__1__61_chany_bottom_out;
wire [0:63] cby_1__1__61_chany_top_out;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__62_ccff_tail;
wire [0:63] cby_1__1__62_chany_bottom_out;
wire [0:63] cby_1__1__62_chany_top_out;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__63_ccff_tail;
wire [0:63] cby_1__1__63_chany_bottom_out;
wire [0:63] cby_1__1__63_chany_top_out;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__64_ccff_tail;
wire [0:63] cby_1__1__64_chany_bottom_out;
wire [0:63] cby_1__1__64_chany_top_out;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__65_ccff_tail;
wire [0:63] cby_1__1__65_chany_bottom_out;
wire [0:63] cby_1__1__65_chany_top_out;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__66_ccff_tail;
wire [0:63] cby_1__1__66_chany_bottom_out;
wire [0:63] cby_1__1__66_chany_top_out;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__67_ccff_tail;
wire [0:63] cby_1__1__67_chany_bottom_out;
wire [0:63] cby_1__1__67_chany_top_out;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__68_ccff_tail;
wire [0:63] cby_1__1__68_chany_bottom_out;
wire [0:63] cby_1__1__68_chany_top_out;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__69_ccff_tail;
wire [0:63] cby_1__1__69_chany_bottom_out;
wire [0:63] cby_1__1__69_chany_top_out;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__6_ccff_tail;
wire [0:63] cby_1__1__6_chany_bottom_out;
wire [0:63] cby_1__1__6_chany_top_out;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__70_ccff_tail;
wire [0:63] cby_1__1__70_chany_bottom_out;
wire [0:63] cby_1__1__70_chany_top_out;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__71_ccff_tail;
wire [0:63] cby_1__1__71_chany_bottom_out;
wire [0:63] cby_1__1__71_chany_top_out;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__72_ccff_tail;
wire [0:63] cby_1__1__72_chany_bottom_out;
wire [0:63] cby_1__1__72_chany_top_out;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__73_ccff_tail;
wire [0:63] cby_1__1__73_chany_bottom_out;
wire [0:63] cby_1__1__73_chany_top_out;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__74_ccff_tail;
wire [0:63] cby_1__1__74_chany_bottom_out;
wire [0:63] cby_1__1__74_chany_top_out;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__75_ccff_tail;
wire [0:63] cby_1__1__75_chany_bottom_out;
wire [0:63] cby_1__1__75_chany_top_out;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__76_ccff_tail;
wire [0:63] cby_1__1__76_chany_bottom_out;
wire [0:63] cby_1__1__76_chany_top_out;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__77_ccff_tail;
wire [0:63] cby_1__1__77_chany_bottom_out;
wire [0:63] cby_1__1__77_chany_top_out;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__78_ccff_tail;
wire [0:63] cby_1__1__78_chany_bottom_out;
wire [0:63] cby_1__1__78_chany_top_out;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__79_ccff_tail;
wire [0:63] cby_1__1__79_chany_bottom_out;
wire [0:63] cby_1__1__79_chany_top_out;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__7_ccff_tail;
wire [0:63] cby_1__1__7_chany_bottom_out;
wire [0:63] cby_1__1__7_chany_top_out;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__80_ccff_tail;
wire [0:63] cby_1__1__80_chany_bottom_out;
wire [0:63] cby_1__1__80_chany_top_out;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__81_ccff_tail;
wire [0:63] cby_1__1__81_chany_bottom_out;
wire [0:63] cby_1__1__81_chany_top_out;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__82_ccff_tail;
wire [0:63] cby_1__1__82_chany_bottom_out;
wire [0:63] cby_1__1__82_chany_top_out;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__83_ccff_tail;
wire [0:63] cby_1__1__83_chany_bottom_out;
wire [0:63] cby_1__1__83_chany_top_out;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__84_ccff_tail;
wire [0:63] cby_1__1__84_chany_bottom_out;
wire [0:63] cby_1__1__84_chany_top_out;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__85_ccff_tail;
wire [0:63] cby_1__1__85_chany_bottom_out;
wire [0:63] cby_1__1__85_chany_top_out;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__86_ccff_tail;
wire [0:63] cby_1__1__86_chany_bottom_out;
wire [0:63] cby_1__1__86_chany_top_out;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__87_ccff_tail;
wire [0:63] cby_1__1__87_chany_bottom_out;
wire [0:63] cby_1__1__87_chany_top_out;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__88_ccff_tail;
wire [0:63] cby_1__1__88_chany_bottom_out;
wire [0:63] cby_1__1__88_chany_top_out;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__89_ccff_tail;
wire [0:63] cby_1__1__89_chany_bottom_out;
wire [0:63] cby_1__1__89_chany_top_out;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__8_ccff_tail;
wire [0:63] cby_1__1__8_chany_bottom_out;
wire [0:63] cby_1__1__8_chany_top_out;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__90_ccff_tail;
wire [0:63] cby_1__1__90_chany_bottom_out;
wire [0:63] cby_1__1__90_chany_top_out;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__91_ccff_tail;
wire [0:63] cby_1__1__91_chany_bottom_out;
wire [0:63] cby_1__1__91_chany_top_out;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__92_ccff_tail;
wire [0:63] cby_1__1__92_chany_bottom_out;
wire [0:63] cby_1__1__92_chany_top_out;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__93_ccff_tail;
wire [0:63] cby_1__1__93_chany_bottom_out;
wire [0:63] cby_1__1__93_chany_top_out;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__94_ccff_tail;
wire [0:63] cby_1__1__94_chany_bottom_out;
wire [0:63] cby_1__1__94_chany_top_out;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__95_ccff_tail;
wire [0:63] cby_1__1__95_chany_bottom_out;
wire [0:63] cby_1__1__95_chany_top_out;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__96_ccff_tail;
wire [0:63] cby_1__1__96_chany_bottom_out;
wire [0:63] cby_1__1__96_chany_top_out;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__97_ccff_tail;
wire [0:63] cby_1__1__97_chany_bottom_out;
wire [0:63] cby_1__1__97_chany_top_out;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__98_ccff_tail;
wire [0:63] cby_1__1__98_chany_bottom_out;
wire [0:63] cby_1__1__98_chany_top_out;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__99_ccff_tail;
wire [0:63] cby_1__1__99_chany_bottom_out;
wire [0:63] cby_1__1__99_chany_top_out;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__9_ccff_tail;
wire [0:63] cby_1__1__9_chany_bottom_out;
wire [0:63] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__0_ccff_tail;
wire [0:63] cby_3__1__0_chany_bottom_out;
wire [0:63] cby_3__1__0_chany_top_out;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__10_ccff_tail;
wire [0:63] cby_3__1__10_chany_bottom_out;
wire [0:63] cby_3__1__10_chany_top_out;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__11_ccff_tail;
wire [0:63] cby_3__1__11_chany_bottom_out;
wire [0:63] cby_3__1__11_chany_top_out;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__12_ccff_tail;
wire [0:63] cby_3__1__12_chany_bottom_out;
wire [0:63] cby_3__1__12_chany_top_out;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__13_ccff_tail;
wire [0:63] cby_3__1__13_chany_bottom_out;
wire [0:63] cby_3__1__13_chany_top_out;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__14_ccff_tail;
wire [0:63] cby_3__1__14_chany_bottom_out;
wire [0:63] cby_3__1__14_chany_top_out;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__15_ccff_tail;
wire [0:63] cby_3__1__15_chany_bottom_out;
wire [0:63] cby_3__1__15_chany_top_out;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__16_ccff_tail;
wire [0:63] cby_3__1__16_chany_bottom_out;
wire [0:63] cby_3__1__16_chany_top_out;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__17_ccff_tail;
wire [0:63] cby_3__1__17_chany_bottom_out;
wire [0:63] cby_3__1__17_chany_top_out;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__1_ccff_tail;
wire [0:63] cby_3__1__1_chany_bottom_out;
wire [0:63] cby_3__1__1_chany_top_out;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__2_ccff_tail;
wire [0:63] cby_3__1__2_chany_bottom_out;
wire [0:63] cby_3__1__2_chany_top_out;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__3_ccff_tail;
wire [0:63] cby_3__1__3_chany_bottom_out;
wire [0:63] cby_3__1__3_chany_top_out;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__4_ccff_tail;
wire [0:63] cby_3__1__4_chany_bottom_out;
wire [0:63] cby_3__1__4_chany_top_out;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__5_ccff_tail;
wire [0:63] cby_3__1__5_chany_bottom_out;
wire [0:63] cby_3__1__5_chany_top_out;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__6_ccff_tail;
wire [0:63] cby_3__1__6_chany_bottom_out;
wire [0:63] cby_3__1__6_chany_top_out;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__7_ccff_tail;
wire [0:63] cby_3__1__7_chany_bottom_out;
wire [0:63] cby_3__1__7_chany_top_out;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__8_ccff_tail;
wire [0:63] cby_3__1__8_chany_bottom_out;
wire [0:63] cby_3__1__8_chany_top_out;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__1__9_ccff_tail;
wire [0:63] cby_3__1__9_chany_bottom_out;
wire [0:63] cby_3__1__9_chany_top_out;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cby_3__2__0_ccff_tail;
wire [0:63] cby_3__2__0_chany_bottom_out;
wire [0:63] cby_3__2__0_chany_top_out;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__10_ccff_tail;
wire [0:63] cby_3__2__10_chany_bottom_out;
wire [0:63] cby_3__2__10_chany_top_out;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__11_ccff_tail;
wire [0:63] cby_3__2__11_chany_bottom_out;
wire [0:63] cby_3__2__11_chany_top_out;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__12_ccff_tail;
wire [0:63] cby_3__2__12_chany_bottom_out;
wire [0:63] cby_3__2__12_chany_top_out;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__13_ccff_tail;
wire [0:63] cby_3__2__13_chany_bottom_out;
wire [0:63] cby_3__2__13_chany_top_out;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__14_ccff_tail;
wire [0:63] cby_3__2__14_chany_bottom_out;
wire [0:63] cby_3__2__14_chany_top_out;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__15_ccff_tail;
wire [0:63] cby_3__2__15_chany_bottom_out;
wire [0:63] cby_3__2__15_chany_top_out;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__16_ccff_tail;
wire [0:63] cby_3__2__16_chany_bottom_out;
wire [0:63] cby_3__2__16_chany_top_out;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__17_ccff_tail;
wire [0:63] cby_3__2__17_chany_bottom_out;
wire [0:63] cby_3__2__17_chany_top_out;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__1_ccff_tail;
wire [0:63] cby_3__2__1_chany_bottom_out;
wire [0:63] cby_3__2__1_chany_top_out;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__2_ccff_tail;
wire [0:63] cby_3__2__2_chany_bottom_out;
wire [0:63] cby_3__2__2_chany_top_out;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__3_ccff_tail;
wire [0:63] cby_3__2__3_chany_bottom_out;
wire [0:63] cby_3__2__3_chany_top_out;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__4_ccff_tail;
wire [0:63] cby_3__2__4_chany_bottom_out;
wire [0:63] cby_3__2__4_chany_top_out;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__5_ccff_tail;
wire [0:63] cby_3__2__5_chany_bottom_out;
wire [0:63] cby_3__2__5_chany_top_out;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__6_ccff_tail;
wire [0:63] cby_3__2__6_chany_bottom_out;
wire [0:63] cby_3__2__6_chany_top_out;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__7_ccff_tail;
wire [0:63] cby_3__2__7_chany_bottom_out;
wire [0:63] cby_3__2__7_chany_top_out;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__8_ccff_tail;
wire [0:63] cby_3__2__8_chany_bottom_out;
wire [0:63] cby_3__2__8_chany_top_out;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_3__2__9_ccff_tail;
wire [0:63] cby_3__2__9_chany_bottom_out;
wire [0:63] cby_3__2__9_chany_top_out;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_;
wire [0:0] cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_;
wire [0:0] cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_;
wire [0:0] cby_4__1__0_ccff_tail;
wire [0:63] cby_4__1__0_chany_bottom_out;
wire [0:63] cby_4__1__0_chany_top_out;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__10_ccff_tail;
wire [0:63] cby_4__1__10_chany_bottom_out;
wire [0:63] cby_4__1__10_chany_top_out;
wire [0:0] cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__11_ccff_tail;
wire [0:63] cby_4__1__11_chany_bottom_out;
wire [0:63] cby_4__1__11_chany_top_out;
wire [0:0] cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__12_ccff_tail;
wire [0:63] cby_4__1__12_chany_bottom_out;
wire [0:63] cby_4__1__12_chany_top_out;
wire [0:0] cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__13_ccff_tail;
wire [0:63] cby_4__1__13_chany_bottom_out;
wire [0:63] cby_4__1__13_chany_top_out;
wire [0:0] cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__14_ccff_tail;
wire [0:63] cby_4__1__14_chany_bottom_out;
wire [0:63] cby_4__1__14_chany_top_out;
wire [0:0] cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__15_ccff_tail;
wire [0:63] cby_4__1__15_chany_bottom_out;
wire [0:63] cby_4__1__15_chany_top_out;
wire [0:0] cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__16_ccff_tail;
wire [0:63] cby_4__1__16_chany_bottom_out;
wire [0:63] cby_4__1__16_chany_top_out;
wire [0:0] cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__17_ccff_tail;
wire [0:63] cby_4__1__17_chany_bottom_out;
wire [0:63] cby_4__1__17_chany_top_out;
wire [0:0] cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__18_ccff_tail;
wire [0:63] cby_4__1__18_chany_bottom_out;
wire [0:63] cby_4__1__18_chany_top_out;
wire [0:0] cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__19_ccff_tail;
wire [0:63] cby_4__1__19_chany_bottom_out;
wire [0:63] cby_4__1__19_chany_top_out;
wire [0:0] cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__1_ccff_tail;
wire [0:63] cby_4__1__1_chany_bottom_out;
wire [0:63] cby_4__1__1_chany_top_out;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__20_ccff_tail;
wire [0:63] cby_4__1__20_chany_bottom_out;
wire [0:63] cby_4__1__20_chany_top_out;
wire [0:0] cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__21_ccff_tail;
wire [0:63] cby_4__1__21_chany_bottom_out;
wire [0:63] cby_4__1__21_chany_top_out;
wire [0:0] cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__22_ccff_tail;
wire [0:63] cby_4__1__22_chany_bottom_out;
wire [0:63] cby_4__1__22_chany_top_out;
wire [0:0] cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__23_ccff_tail;
wire [0:63] cby_4__1__23_chany_bottom_out;
wire [0:63] cby_4__1__23_chany_top_out;
wire [0:0] cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__24_ccff_tail;
wire [0:63] cby_4__1__24_chany_bottom_out;
wire [0:63] cby_4__1__24_chany_top_out;
wire [0:0] cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__25_ccff_tail;
wire [0:63] cby_4__1__25_chany_bottom_out;
wire [0:63] cby_4__1__25_chany_top_out;
wire [0:0] cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__26_ccff_tail;
wire [0:63] cby_4__1__26_chany_bottom_out;
wire [0:63] cby_4__1__26_chany_top_out;
wire [0:0] cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__27_ccff_tail;
wire [0:63] cby_4__1__27_chany_bottom_out;
wire [0:63] cby_4__1__27_chany_top_out;
wire [0:0] cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__28_ccff_tail;
wire [0:63] cby_4__1__28_chany_bottom_out;
wire [0:63] cby_4__1__28_chany_top_out;
wire [0:0] cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__29_ccff_tail;
wire [0:63] cby_4__1__29_chany_bottom_out;
wire [0:63] cby_4__1__29_chany_top_out;
wire [0:0] cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__2_ccff_tail;
wire [0:63] cby_4__1__2_chany_bottom_out;
wire [0:63] cby_4__1__2_chany_top_out;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:63] cby_4__1__30_chany_bottom_out;
wire [0:63] cby_4__1__30_chany_top_out;
wire [0:0] cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__31_ccff_tail;
wire [0:63] cby_4__1__31_chany_bottom_out;
wire [0:63] cby_4__1__31_chany_top_out;
wire [0:0] cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__32_ccff_tail;
wire [0:63] cby_4__1__32_chany_bottom_out;
wire [0:63] cby_4__1__32_chany_top_out;
wire [0:0] cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__33_ccff_tail;
wire [0:63] cby_4__1__33_chany_bottom_out;
wire [0:63] cby_4__1__33_chany_top_out;
wire [0:0] cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__34_ccff_tail;
wire [0:63] cby_4__1__34_chany_bottom_out;
wire [0:63] cby_4__1__34_chany_top_out;
wire [0:0] cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__35_ccff_tail;
wire [0:63] cby_4__1__35_chany_bottom_out;
wire [0:63] cby_4__1__35_chany_top_out;
wire [0:0] cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__3_ccff_tail;
wire [0:63] cby_4__1__3_chany_bottom_out;
wire [0:63] cby_4__1__3_chany_top_out;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__4_ccff_tail;
wire [0:63] cby_4__1__4_chany_bottom_out;
wire [0:63] cby_4__1__4_chany_top_out;
wire [0:0] cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__5_ccff_tail;
wire [0:63] cby_4__1__5_chany_bottom_out;
wire [0:63] cby_4__1__5_chany_top_out;
wire [0:0] cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__6_ccff_tail;
wire [0:63] cby_4__1__6_chany_bottom_out;
wire [0:63] cby_4__1__6_chany_top_out;
wire [0:0] cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__7_ccff_tail;
wire [0:63] cby_4__1__7_chany_bottom_out;
wire [0:63] cby_4__1__7_chany_top_out;
wire [0:0] cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__8_ccff_tail;
wire [0:63] cby_4__1__8_chany_bottom_out;
wire [0:63] cby_4__1__8_chany_top_out;
wire [0:0] cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_4__1__9_ccff_tail;
wire [0:63] cby_4__1__9_chany_bottom_out;
wire [0:63] cby_4__1__9_chany_top_out;
wire [0:0] cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_100_out;
wire [0:0] direct_interc_101_out;
wire [0:0] direct_interc_102_out;
wire [0:0] direct_interc_103_out;
wire [0:0] direct_interc_104_out;
wire [0:0] direct_interc_105_out;
wire [0:0] direct_interc_106_out;
wire [0:0] direct_interc_107_out;
wire [0:0] direct_interc_108_out;
wire [0:0] direct_interc_109_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_110_out;
wire [0:0] direct_interc_111_out;
wire [0:0] direct_interc_112_out;
wire [0:0] direct_interc_113_out;
wire [0:0] direct_interc_114_out;
wire [0:0] direct_interc_115_out;
wire [0:0] direct_interc_116_out;
wire [0:0] direct_interc_117_out;
wire [0:0] direct_interc_118_out;
wire [0:0] direct_interc_119_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_120_out;
wire [0:0] direct_interc_121_out;
wire [0:0] direct_interc_122_out;
wire [0:0] direct_interc_123_out;
wire [0:0] direct_interc_124_out;
wire [0:0] direct_interc_125_out;
wire [0:0] direct_interc_126_out;
wire [0:0] direct_interc_127_out;
wire [0:0] direct_interc_128_out;
wire [0:0] direct_interc_129_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_130_out;
wire [0:0] direct_interc_131_out;
wire [0:0] direct_interc_132_out;
wire [0:0] direct_interc_133_out;
wire [0:0] direct_interc_134_out;
wire [0:0] direct_interc_135_out;
wire [0:0] direct_interc_136_out;
wire [0:0] direct_interc_137_out;
wire [0:0] direct_interc_138_out;
wire [0:0] direct_interc_139_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_140_out;
wire [0:0] direct_interc_141_out;
wire [0:0] direct_interc_142_out;
wire [0:0] direct_interc_143_out;
wire [0:0] direct_interc_144_out;
wire [0:0] direct_interc_145_out;
wire [0:0] direct_interc_146_out;
wire [0:0] direct_interc_147_out;
wire [0:0] direct_interc_148_out;
wire [0:0] direct_interc_149_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_150_out;
wire [0:0] direct_interc_151_out;
wire [0:0] direct_interc_152_out;
wire [0:0] direct_interc_153_out;
wire [0:0] direct_interc_154_out;
wire [0:0] direct_interc_155_out;
wire [0:0] direct_interc_156_out;
wire [0:0] direct_interc_157_out;
wire [0:0] direct_interc_158_out;
wire [0:0] direct_interc_159_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_160_out;
wire [0:0] direct_interc_161_out;
wire [0:0] direct_interc_162_out;
wire [0:0] direct_interc_163_out;
wire [0:0] direct_interc_164_out;
wire [0:0] direct_interc_165_out;
wire [0:0] direct_interc_166_out;
wire [0:0] direct_interc_167_out;
wire [0:0] direct_interc_168_out;
wire [0:0] direct_interc_169_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_170_out;
wire [0:0] direct_interc_171_out;
wire [0:0] direct_interc_172_out;
wire [0:0] direct_interc_173_out;
wire [0:0] direct_interc_174_out;
wire [0:0] direct_interc_175_out;
wire [0:0] direct_interc_176_out;
wire [0:0] direct_interc_177_out;
wire [0:0] direct_interc_178_out;
wire [0:0] direct_interc_179_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_180_out;
wire [0:0] direct_interc_181_out;
wire [0:0] direct_interc_182_out;
wire [0:0] direct_interc_183_out;
wire [0:0] direct_interc_184_out;
wire [0:0] direct_interc_185_out;
wire [0:0] direct_interc_186_out;
wire [0:0] direct_interc_187_out;
wire [0:0] direct_interc_188_out;
wire [0:0] direct_interc_189_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_190_out;
wire [0:0] direct_interc_191_out;
wire [0:0] direct_interc_192_out;
wire [0:0] direct_interc_193_out;
wire [0:0] direct_interc_194_out;
wire [0:0] direct_interc_195_out;
wire [0:0] direct_interc_196_out;
wire [0:0] direct_interc_197_out;
wire [0:0] direct_interc_198_out;
wire [0:0] direct_interc_199_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_200_out;
wire [0:0] direct_interc_201_out;
wire [0:0] direct_interc_202_out;
wire [0:0] direct_interc_203_out;
wire [0:0] direct_interc_204_out;
wire [0:0] direct_interc_205_out;
wire [0:0] direct_interc_206_out;
wire [0:0] direct_interc_207_out;
wire [0:0] direct_interc_208_out;
wire [0:0] direct_interc_209_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_210_out;
wire [0:0] direct_interc_211_out;
wire [0:0] direct_interc_212_out;
wire [0:0] direct_interc_213_out;
wire [0:0] direct_interc_214_out;
wire [0:0] direct_interc_215_out;
wire [0:0] direct_interc_216_out;
wire [0:0] direct_interc_217_out;
wire [0:0] direct_interc_218_out;
wire [0:0] direct_interc_219_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_220_out;
wire [0:0] direct_interc_221_out;
wire [0:0] direct_interc_222_out;
wire [0:0] direct_interc_223_out;
wire [0:0] direct_interc_224_out;
wire [0:0] direct_interc_225_out;
wire [0:0] direct_interc_226_out;
wire [0:0] direct_interc_227_out;
wire [0:0] direct_interc_228_out;
wire [0:0] direct_interc_229_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_230_out;
wire [0:0] direct_interc_231_out;
wire [0:0] direct_interc_232_out;
wire [0:0] direct_interc_233_out;
wire [0:0] direct_interc_234_out;
wire [0:0] direct_interc_235_out;
wire [0:0] direct_interc_236_out;
wire [0:0] direct_interc_237_out;
wire [0:0] direct_interc_238_out;
wire [0:0] direct_interc_239_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_240_out;
wire [0:0] direct_interc_241_out;
wire [0:0] direct_interc_242_out;
wire [0:0] direct_interc_243_out;
wire [0:0] direct_interc_244_out;
wire [0:0] direct_interc_245_out;
wire [0:0] direct_interc_246_out;
wire [0:0] direct_interc_247_out;
wire [0:0] direct_interc_248_out;
wire [0:0] direct_interc_249_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_250_out;
wire [0:0] direct_interc_251_out;
wire [0:0] direct_interc_252_out;
wire [0:0] direct_interc_253_out;
wire [0:0] direct_interc_254_out;
wire [0:0] direct_interc_255_out;
wire [0:0] direct_interc_256_out;
wire [0:0] direct_interc_257_out;
wire [0:0] direct_interc_258_out;
wire [0:0] direct_interc_259_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_260_out;
wire [0:0] direct_interc_261_out;
wire [0:0] direct_interc_262_out;
wire [0:0] direct_interc_263_out;
wire [0:0] direct_interc_264_out;
wire [0:0] direct_interc_265_out;
wire [0:0] direct_interc_266_out;
wire [0:0] direct_interc_267_out;
wire [0:0] direct_interc_268_out;
wire [0:0] direct_interc_269_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_270_out;
wire [0:0] direct_interc_271_out;
wire [0:0] direct_interc_272_out;
wire [0:0] direct_interc_273_out;
wire [0:0] direct_interc_274_out;
wire [0:0] direct_interc_275_out;
wire [0:0] direct_interc_276_out;
wire [0:0] direct_interc_277_out;
wire [0:0] direct_interc_278_out;
wire [0:0] direct_interc_279_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_280_out;
wire [0:0] direct_interc_281_out;
wire [0:0] direct_interc_282_out;
wire [0:0] direct_interc_283_out;
wire [0:0] direct_interc_284_out;
wire [0:0] direct_interc_285_out;
wire [0:0] direct_interc_286_out;
wire [0:0] direct_interc_287_out;
wire [0:0] direct_interc_288_out;
wire [0:0] direct_interc_289_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_290_out;
wire [0:0] direct_interc_291_out;
wire [0:0] direct_interc_292_out;
wire [0:0] direct_interc_293_out;
wire [0:0] direct_interc_294_out;
wire [0:0] direct_interc_295_out;
wire [0:0] direct_interc_296_out;
wire [0:0] direct_interc_297_out;
wire [0:0] direct_interc_298_out;
wire [0:0] direct_interc_299_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_300_out;
wire [0:0] direct_interc_301_out;
wire [0:0] direct_interc_302_out;
wire [0:0] direct_interc_303_out;
wire [0:0] direct_interc_304_out;
wire [0:0] direct_interc_305_out;
wire [0:0] direct_interc_306_out;
wire [0:0] direct_interc_307_out;
wire [0:0] direct_interc_308_out;
wire [0:0] direct_interc_309_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_310_out;
wire [0:0] direct_interc_311_out;
wire [0:0] direct_interc_312_out;
wire [0:0] direct_interc_313_out;
wire [0:0] direct_interc_314_out;
wire [0:0] direct_interc_315_out;
wire [0:0] direct_interc_316_out;
wire [0:0] direct_interc_317_out;
wire [0:0] direct_interc_318_out;
wire [0:0] direct_interc_319_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_320_out;
wire [0:0] direct_interc_321_out;
wire [0:0] direct_interc_322_out;
wire [0:0] direct_interc_323_out;
wire [0:0] direct_interc_324_out;
wire [0:0] direct_interc_325_out;
wire [0:0] direct_interc_326_out;
wire [0:0] direct_interc_327_out;
wire [0:0] direct_interc_328_out;
wire [0:0] direct_interc_329_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_330_out;
wire [0:0] direct_interc_331_out;
wire [0:0] direct_interc_332_out;
wire [0:0] direct_interc_333_out;
wire [0:0] direct_interc_334_out;
wire [0:0] direct_interc_335_out;
wire [0:0] direct_interc_336_out;
wire [0:0] direct_interc_337_out;
wire [0:0] direct_interc_338_out;
wire [0:0] direct_interc_339_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_340_out;
wire [0:0] direct_interc_341_out;
wire [0:0] direct_interc_342_out;
wire [0:0] direct_interc_343_out;
wire [0:0] direct_interc_344_out;
wire [0:0] direct_interc_345_out;
wire [0:0] direct_interc_346_out;
wire [0:0] direct_interc_347_out;
wire [0:0] direct_interc_348_out;
wire [0:0] direct_interc_349_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_350_out;
wire [0:0] direct_interc_351_out;
wire [0:0] direct_interc_352_out;
wire [0:0] direct_interc_353_out;
wire [0:0] direct_interc_354_out;
wire [0:0] direct_interc_355_out;
wire [0:0] direct_interc_356_out;
wire [0:0] direct_interc_357_out;
wire [0:0] direct_interc_358_out;
wire [0:0] direct_interc_359_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_360_out;
wire [0:0] direct_interc_361_out;
wire [0:0] direct_interc_362_out;
wire [0:0] direct_interc_363_out;
wire [0:0] direct_interc_364_out;
wire [0:0] direct_interc_365_out;
wire [0:0] direct_interc_366_out;
wire [0:0] direct_interc_367_out;
wire [0:0] direct_interc_368_out;
wire [0:0] direct_interc_369_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_370_out;
wire [0:0] direct_interc_371_out;
wire [0:0] direct_interc_372_out;
wire [0:0] direct_interc_373_out;
wire [0:0] direct_interc_374_out;
wire [0:0] direct_interc_375_out;
wire [0:0] direct_interc_376_out;
wire [0:0] direct_interc_377_out;
wire [0:0] direct_interc_378_out;
wire [0:0] direct_interc_379_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_380_out;
wire [0:0] direct_interc_381_out;
wire [0:0] direct_interc_382_out;
wire [0:0] direct_interc_383_out;
wire [0:0] direct_interc_384_out;
wire [0:0] direct_interc_385_out;
wire [0:0] direct_interc_386_out;
wire [0:0] direct_interc_387_out;
wire [0:0] direct_interc_388_out;
wire [0:0] direct_interc_389_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_390_out;
wire [0:0] direct_interc_391_out;
wire [0:0] direct_interc_392_out;
wire [0:0] direct_interc_393_out;
wire [0:0] direct_interc_394_out;
wire [0:0] direct_interc_395_out;
wire [0:0] direct_interc_396_out;
wire [0:0] direct_interc_397_out;
wire [0:0] direct_interc_398_out;
wire [0:0] direct_interc_399_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_400_out;
wire [0:0] direct_interc_401_out;
wire [0:0] direct_interc_402_out;
wire [0:0] direct_interc_403_out;
wire [0:0] direct_interc_404_out;
wire [0:0] direct_interc_405_out;
wire [0:0] direct_interc_406_out;
wire [0:0] direct_interc_407_out;
wire [0:0] direct_interc_408_out;
wire [0:0] direct_interc_409_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_410_out;
wire [0:0] direct_interc_411_out;
wire [0:0] direct_interc_412_out;
wire [0:0] direct_interc_413_out;
wire [0:0] direct_interc_414_out;
wire [0:0] direct_interc_415_out;
wire [0:0] direct_interc_416_out;
wire [0:0] direct_interc_417_out;
wire [0:0] direct_interc_418_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_44_out;
wire [0:0] direct_interc_45_out;
wire [0:0] direct_interc_46_out;
wire [0:0] direct_interc_47_out;
wire [0:0] direct_interc_48_out;
wire [0:0] direct_interc_49_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_50_out;
wire [0:0] direct_interc_51_out;
wire [0:0] direct_interc_52_out;
wire [0:0] direct_interc_53_out;
wire [0:0] direct_interc_54_out;
wire [0:0] direct_interc_55_out;
wire [0:0] direct_interc_56_out;
wire [0:0] direct_interc_57_out;
wire [0:0] direct_interc_58_out;
wire [0:0] direct_interc_59_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_60_out;
wire [0:0] direct_interc_61_out;
wire [0:0] direct_interc_62_out;
wire [0:0] direct_interc_63_out;
wire [0:0] direct_interc_64_out;
wire [0:0] direct_interc_65_out;
wire [0:0] direct_interc_66_out;
wire [0:0] direct_interc_67_out;
wire [0:0] direct_interc_68_out;
wire [0:0] direct_interc_69_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_70_out;
wire [0:0] direct_interc_71_out;
wire [0:0] direct_interc_72_out;
wire [0:0] direct_interc_73_out;
wire [0:0] direct_interc_74_out;
wire [0:0] direct_interc_75_out;
wire [0:0] direct_interc_76_out;
wire [0:0] direct_interc_77_out;
wire [0:0] direct_interc_78_out;
wire [0:0] direct_interc_79_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_80_out;
wire [0:0] direct_interc_81_out;
wire [0:0] direct_interc_82_out;
wire [0:0] direct_interc_83_out;
wire [0:0] direct_interc_84_out;
wire [0:0] direct_interc_85_out;
wire [0:0] direct_interc_86_out;
wire [0:0] direct_interc_87_out;
wire [0:0] direct_interc_88_out;
wire [0:0] direct_interc_89_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_90_out;
wire [0:0] direct_interc_91_out;
wire [0:0] direct_interc_92_out;
wire [0:0] direct_interc_93_out;
wire [0:0] direct_interc_94_out;
wire [0:0] direct_interc_95_out;
wire [0:0] direct_interc_96_out;
wire [0:0] direct_interc_97_out;
wire [0:0] direct_interc_98_out;
wire [0:0] direct_interc_99_out;
wire [0:0] direct_interc_9_out;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_100_ccff_tail;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_101_ccff_tail;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_102_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_102_ccff_tail;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_103_ccff_tail;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_104_ccff_tail;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_105_ccff_tail;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_106_ccff_tail;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_107_ccff_tail;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_108_ccff_tail;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_109_ccff_tail;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_10__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_110_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_110_ccff_tail;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_111_ccff_tail;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_112_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_112_ccff_tail;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_113_ccff_tail;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_114_ccff_tail;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_115_ccff_tail;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_116_ccff_tail;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_117_ccff_tail;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_118_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_118_ccff_tail;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_119_ccff_tail;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_120_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_120_ccff_tail;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_121_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_121_ccff_tail;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_122_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_122_ccff_tail;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_123_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_123_ccff_tail;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_124_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_124_ccff_tail;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_125_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_125_ccff_tail;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_126_ccff_tail;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_127_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_127_ccff_tail;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_128_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_128_ccff_tail;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_129_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_129_ccff_tail;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_12__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_130_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_130_ccff_tail;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_131_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_131_ccff_tail;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_132_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_132_ccff_tail;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_133_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_133_ccff_tail;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_134_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_134_ccff_tail;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_135_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_135_ccff_tail;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_136_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_136_ccff_tail;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_137_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_137_ccff_tail;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_138_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_138_ccff_tail;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_139_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_139_ccff_tail;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_13__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_13__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_140_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_140_ccff_tail;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_141_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_141_ccff_tail;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_142_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_142_ccff_tail;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_143_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_143_ccff_tail;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_144_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_144_ccff_tail;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_145_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_145_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_145_ccff_tail;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_146_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_146_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_146_ccff_tail;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_147_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_147_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_147_ccff_tail;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_148_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_148_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_148_ccff_tail;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_149_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_149_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_149_ccff_tail;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_14__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_14__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_14__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_150_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_150_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_150_ccff_tail;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_151_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_151_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_151_ccff_tail;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_152_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_152_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_152_ccff_tail;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_153_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_153_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_153_ccff_tail;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_154_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_154_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_154_ccff_tail;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_155_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_155_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_155_ccff_tail;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_156_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_156_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_156_ccff_tail;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_157_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_157_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_157_ccff_tail;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_158_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_158_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_158_ccff_tail;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_159_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_159_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_159_ccff_tail;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_160_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_160_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_160_ccff_tail;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_161_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_161_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_161_ccff_tail;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_162_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_162_ccff_tail;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_163_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_163_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_163_ccff_tail;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_164_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_164_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_164_ccff_tail;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_165_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_165_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_165_ccff_tail;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_166_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_166_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_166_ccff_tail;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_167_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_167_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_167_ccff_tail;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_168_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_168_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_168_ccff_tail;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_169_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_169_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_169_ccff_tail;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_170_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_170_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_170_ccff_tail;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_171_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_171_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_171_ccff_tail;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_172_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_172_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_172_ccff_tail;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_173_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_173_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_173_ccff_tail;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_174_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_174_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_174_ccff_tail;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_175_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_175_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_175_ccff_tail;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_176_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_176_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_176_ccff_tail;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_177_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_177_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_177_ccff_tail;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_178_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_178_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_178_ccff_tail;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_179_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_179_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_179_ccff_tail;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_180_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_180_ccff_tail;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_181_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_181_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_181_ccff_tail;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_182_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_182_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_182_ccff_tail;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_183_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_183_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_183_ccff_tail;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_184_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_184_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_184_ccff_tail;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_185_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_185_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_185_ccff_tail;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_186_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_186_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_186_ccff_tail;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_187_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_187_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_187_ccff_tail;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_188_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_188_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_188_ccff_tail;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_189_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_189_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_189_ccff_tail;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_190_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_190_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_190_ccff_tail;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_191_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_191_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_191_ccff_tail;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_192_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_192_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_192_ccff_tail;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_193_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_193_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_193_ccff_tail;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_194_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_194_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_194_ccff_tail;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_195_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_195_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_195_ccff_tail;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_196_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_196_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_196_ccff_tail;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_197_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_197_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_197_ccff_tail;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_198_ccff_tail;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_199_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_199_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_199_ccff_tail;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_1__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__18__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_200_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_200_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_200_ccff_tail;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_201_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_201_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_201_ccff_tail;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_202_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_202_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_202_ccff_tail;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_203_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_203_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_203_ccff_tail;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_204_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_204_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_204_ccff_tail;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_205_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_205_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_205_ccff_tail;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_206_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_206_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_206_ccff_tail;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_207_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_207_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_207_ccff_tail;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_208_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_208_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_208_ccff_tail;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_209_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_209_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_209_ccff_tail;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_210_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_210_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_210_ccff_tail;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_211_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_211_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_211_ccff_tail;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_212_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_212_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_212_ccff_tail;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_213_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_213_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_213_ccff_tail;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_214_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_214_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_214_ccff_tail;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_215_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_215_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_215_ccff_tail;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_22_ccff_tail;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_23_ccff_tail;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_24_ccff_tail;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_25_ccff_tail;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_26_ccff_tail;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_27_ccff_tail;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_28_ccff_tail;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_29_ccff_tail;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_2__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_30_ccff_tail;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_31_ccff_tail;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_32_ccff_tail;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_33_ccff_tail;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_35_ccff_tail;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_36_ccff_tail;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_37_ccff_tail;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_38_ccff_tail;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_39_ccff_tail;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_3__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_40_ccff_tail;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_41_ccff_tail;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_42_ccff_tail;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_43_ccff_tail;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_44_ccff_tail;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_45_ccff_tail;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_46_ccff_tail;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_47_ccff_tail;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_48_ccff_tail;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_49_ccff_tail;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_50_ccff_tail;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_51_ccff_tail;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_52_ccff_tail;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_53_ccff_tail;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_54_ccff_tail;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_55_ccff_tail;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_56_ccff_tail;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_57_ccff_tail;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_59_ccff_tail;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_5__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_60_ccff_tail;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_62_ccff_tail;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_63_ccff_tail;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_64_ccff_tail;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_65_ccff_tail;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_66_ccff_tail;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_67_ccff_tail;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_68_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_68_ccff_tail;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_69_ccff_tail;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_6__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_70_ccff_tail;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_71_ccff_tail;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_72_ccff_tail;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_73_ccff_tail;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_74_ccff_tail;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_75_ccff_tail;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_76_ccff_tail;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_77_ccff_tail;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_78_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_78_ccff_tail;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_79_ccff_tail;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_7__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_80_ccff_tail;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_81_ccff_tail;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_82_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_82_ccff_tail;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_83_ccff_tail;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_84_ccff_tail;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_85_ccff_tail;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_86_ccff_tail;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_87_ccff_tail;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_88_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_88_ccff_tail;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_89_ccff_tail;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_8__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_90_ccff_tail;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_91_ccff_tail;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_92_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_92_ccff_tail;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_93_ccff_tail;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_94_ccff_tail;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_95_ccff_tail;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_96_ccff_tail;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_97_ccff_tail;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_98_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_98_ccff_tail;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_99_ccff_tail;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_9__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_ccff_tail;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_ccff_tail;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_ccff_tail;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_ccff_tail;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_ccff_tail;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_ccff_tail;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_ccff_tail;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_ccff_tail;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_0_ccff_tail;
wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_10_ccff_tail;
wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_11_ccff_tail;
wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_12_ccff_tail;
wire [0:0] grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_13_ccff_tail;
wire [0:0] grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_14_ccff_tail;
wire [0:0] grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_15_ccff_tail;
wire [0:0] grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_16_ccff_tail;
wire [0:0] grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_17_ccff_tail;
wire [0:0] grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_1_ccff_tail;
wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_2_ccff_tail;
wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_3_ccff_tail;
wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_4_ccff_tail;
wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_5_ccff_tail;
wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_6_ccff_tail;
wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_7_ccff_tail;
wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_8_ccff_tail;
wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_9_ccff_tail;
wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_0_ccff_tail;
wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_10_ccff_tail;
wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_11_ccff_tail;
wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_12_ccff_tail;
wire [0:0] grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_13_ccff_tail;
wire [0:0] grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_14_ccff_tail;
wire [0:0] grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_15_ccff_tail;
wire [0:0] grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_16_ccff_tail;
wire [0:0] grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_17_ccff_tail;
wire [0:0] grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_1_ccff_tail;
wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_2_ccff_tail;
wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_3_ccff_tail;
wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_4_ccff_tail;
wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_5_ccff_tail;
wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_6_ccff_tail;
wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_7_ccff_tail;
wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_8_ccff_tail;
wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_9_ccff_tail;
wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_0_ccff_tail;
wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_10_ccff_tail;
wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_11_ccff_tail;
wire [0:0] grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_12_ccff_tail;
wire [0:0] grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_13_ccff_tail;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_1_ccff_tail;
wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_2_ccff_tail;
wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_3_ccff_tail;
wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_4_ccff_tail;
wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_5_ccff_tail;
wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_6_ccff_tail;
wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_7_ccff_tail;
wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_8_ccff_tail;
wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_9_ccff_tail;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__13__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__15__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__17__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__13__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__15__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__17__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower;
wire [0:0] grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper;
wire [0:0] grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower;
wire [0:0] grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper;
wire [0:0] grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_lower;
wire [0:0] grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_upper;
wire [0:0] grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_lower;
wire [0:0] grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_upper;
wire [0:0] grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_lower;
wire [0:0] grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_upper;
wire [0:0] grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_lower;
wire [0:0] grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_upper;
wire [0:0] grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_lower;
wire [0:0] grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_upper;
wire [0:0] grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_lower;
wire [0:0] grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_upper;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:63] sb_0__0__0_chanx_right_out;
wire [0:63] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__18__0_ccff_tail;
wire [0:63] sb_0__18__0_chanx_right_out;
wire [0:63] sb_0__18__0_chany_bottom_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:63] sb_0__1__0_chanx_right_out;
wire [0:63] sb_0__1__0_chany_bottom_out;
wire [0:63] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__10_ccff_tail;
wire [0:63] sb_0__1__10_chanx_right_out;
wire [0:63] sb_0__1__10_chany_bottom_out;
wire [0:63] sb_0__1__10_chany_top_out;
wire [0:63] sb_0__1__11_chanx_right_out;
wire [0:63] sb_0__1__11_chany_bottom_out;
wire [0:63] sb_0__1__11_chany_top_out;
wire [0:0] sb_0__1__12_ccff_tail;
wire [0:63] sb_0__1__12_chanx_right_out;
wire [0:63] sb_0__1__12_chany_bottom_out;
wire [0:63] sb_0__1__12_chany_top_out;
wire [0:0] sb_0__1__13_ccff_tail;
wire [0:63] sb_0__1__13_chanx_right_out;
wire [0:63] sb_0__1__13_chany_bottom_out;
wire [0:63] sb_0__1__13_chany_top_out;
wire [0:0] sb_0__1__14_ccff_tail;
wire [0:63] sb_0__1__14_chanx_right_out;
wire [0:63] sb_0__1__14_chany_bottom_out;
wire [0:63] sb_0__1__14_chany_top_out;
wire [0:0] sb_0__1__15_ccff_tail;
wire [0:63] sb_0__1__15_chanx_right_out;
wire [0:63] sb_0__1__15_chany_bottom_out;
wire [0:63] sb_0__1__15_chany_top_out;
wire [0:0] sb_0__1__16_ccff_tail;
wire [0:63] sb_0__1__16_chanx_right_out;
wire [0:63] sb_0__1__16_chany_bottom_out;
wire [0:63] sb_0__1__16_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:63] sb_0__1__1_chanx_right_out;
wire [0:63] sb_0__1__1_chany_bottom_out;
wire [0:63] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__1__2_ccff_tail;
wire [0:63] sb_0__1__2_chanx_right_out;
wire [0:63] sb_0__1__2_chany_bottom_out;
wire [0:63] sb_0__1__2_chany_top_out;
wire [0:0] sb_0__1__3_ccff_tail;
wire [0:63] sb_0__1__3_chanx_right_out;
wire [0:63] sb_0__1__3_chany_bottom_out;
wire [0:63] sb_0__1__3_chany_top_out;
wire [0:0] sb_0__1__4_ccff_tail;
wire [0:63] sb_0__1__4_chanx_right_out;
wire [0:63] sb_0__1__4_chany_bottom_out;
wire [0:63] sb_0__1__4_chany_top_out;
wire [0:0] sb_0__1__5_ccff_tail;
wire [0:63] sb_0__1__5_chanx_right_out;
wire [0:63] sb_0__1__5_chany_bottom_out;
wire [0:63] sb_0__1__5_chany_top_out;
wire [0:0] sb_0__1__6_ccff_tail;
wire [0:63] sb_0__1__6_chanx_right_out;
wire [0:63] sb_0__1__6_chany_bottom_out;
wire [0:63] sb_0__1__6_chany_top_out;
wire [0:0] sb_0__1__7_ccff_tail;
wire [0:63] sb_0__1__7_chanx_right_out;
wire [0:63] sb_0__1__7_chany_bottom_out;
wire [0:63] sb_0__1__7_chany_top_out;
wire [0:0] sb_0__1__8_ccff_tail;
wire [0:63] sb_0__1__8_chanx_right_out;
wire [0:63] sb_0__1__8_chany_bottom_out;
wire [0:63] sb_0__1__8_chany_top_out;
wire [0:0] sb_0__1__9_ccff_tail;
wire [0:63] sb_0__1__9_chanx_right_out;
wire [0:63] sb_0__1__9_chany_bottom_out;
wire [0:63] sb_0__1__9_chany_top_out;
wire [0:0] sb_14__0__0_ccff_tail;
wire [0:63] sb_14__0__0_chanx_left_out;
wire [0:63] sb_14__0__0_chany_top_out;
wire [0:0] sb_14__18__0_ccff_tail;
wire [0:63] sb_14__18__0_chanx_left_out;
wire [0:63] sb_14__18__0_chany_bottom_out;
wire [0:0] sb_14__1__0_ccff_tail;
wire [0:63] sb_14__1__0_chanx_left_out;
wire [0:63] sb_14__1__0_chany_bottom_out;
wire [0:63] sb_14__1__0_chany_top_out;
wire [0:0] sb_14__1__10_ccff_tail;
wire [0:63] sb_14__1__10_chanx_left_out;
wire [0:63] sb_14__1__10_chany_bottom_out;
wire [0:63] sb_14__1__10_chany_top_out;
wire [0:0] sb_14__1__11_ccff_tail;
wire [0:63] sb_14__1__11_chanx_left_out;
wire [0:63] sb_14__1__11_chany_bottom_out;
wire [0:63] sb_14__1__11_chany_top_out;
wire [0:0] sb_14__1__12_ccff_tail;
wire [0:63] sb_14__1__12_chanx_left_out;
wire [0:63] sb_14__1__12_chany_bottom_out;
wire [0:63] sb_14__1__12_chany_top_out;
wire [0:0] sb_14__1__13_ccff_tail;
wire [0:63] sb_14__1__13_chanx_left_out;
wire [0:63] sb_14__1__13_chany_bottom_out;
wire [0:63] sb_14__1__13_chany_top_out;
wire [0:0] sb_14__1__14_ccff_tail;
wire [0:63] sb_14__1__14_chanx_left_out;
wire [0:63] sb_14__1__14_chany_bottom_out;
wire [0:63] sb_14__1__14_chany_top_out;
wire [0:0] sb_14__1__15_ccff_tail;
wire [0:63] sb_14__1__15_chanx_left_out;
wire [0:63] sb_14__1__15_chany_bottom_out;
wire [0:63] sb_14__1__15_chany_top_out;
wire [0:0] sb_14__1__16_ccff_tail;
wire [0:63] sb_14__1__16_chanx_left_out;
wire [0:63] sb_14__1__16_chany_bottom_out;
wire [0:63] sb_14__1__16_chany_top_out;
wire [0:0] sb_14__1__1_ccff_tail;
wire [0:63] sb_14__1__1_chanx_left_out;
wire [0:63] sb_14__1__1_chany_bottom_out;
wire [0:63] sb_14__1__1_chany_top_out;
wire [0:0] sb_14__1__2_ccff_tail;
wire [0:63] sb_14__1__2_chanx_left_out;
wire [0:63] sb_14__1__2_chany_bottom_out;
wire [0:63] sb_14__1__2_chany_top_out;
wire [0:0] sb_14__1__3_ccff_tail;
wire [0:63] sb_14__1__3_chanx_left_out;
wire [0:63] sb_14__1__3_chany_bottom_out;
wire [0:63] sb_14__1__3_chany_top_out;
wire [0:0] sb_14__1__4_ccff_tail;
wire [0:63] sb_14__1__4_chanx_left_out;
wire [0:63] sb_14__1__4_chany_bottom_out;
wire [0:63] sb_14__1__4_chany_top_out;
wire [0:0] sb_14__1__5_ccff_tail;
wire [0:63] sb_14__1__5_chanx_left_out;
wire [0:63] sb_14__1__5_chany_bottom_out;
wire [0:63] sb_14__1__5_chany_top_out;
wire [0:0] sb_14__1__6_ccff_tail;
wire [0:63] sb_14__1__6_chanx_left_out;
wire [0:63] sb_14__1__6_chany_bottom_out;
wire [0:63] sb_14__1__6_chany_top_out;
wire [0:0] sb_14__1__7_ccff_tail;
wire [0:63] sb_14__1__7_chanx_left_out;
wire [0:63] sb_14__1__7_chany_bottom_out;
wire [0:63] sb_14__1__7_chany_top_out;
wire [0:0] sb_14__1__8_ccff_tail;
wire [0:63] sb_14__1__8_chanx_left_out;
wire [0:63] sb_14__1__8_chany_bottom_out;
wire [0:63] sb_14__1__8_chany_top_out;
wire [0:0] sb_14__1__9_ccff_tail;
wire [0:63] sb_14__1__9_chanx_left_out;
wire [0:63] sb_14__1__9_chany_bottom_out;
wire [0:63] sb_14__1__9_chany_top_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:63] sb_1__0__0_chanx_left_out;
wire [0:63] sb_1__0__0_chanx_right_out;
wire [0:63] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:63] sb_1__0__1_chanx_left_out;
wire [0:63] sb_1__0__1_chanx_right_out;
wire [0:63] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:63] sb_1__0__2_chanx_left_out;
wire [0:63] sb_1__0__2_chanx_right_out;
wire [0:63] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:63] sb_1__0__3_chanx_left_out;
wire [0:63] sb_1__0__3_chanx_right_out;
wire [0:63] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:63] sb_1__0__4_chanx_left_out;
wire [0:63] sb_1__0__4_chanx_right_out;
wire [0:63] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__0__5_ccff_tail;
wire [0:63] sb_1__0__5_chanx_left_out;
wire [0:63] sb_1__0__5_chanx_right_out;
wire [0:63] sb_1__0__5_chany_top_out;
wire [0:0] sb_1__0__6_ccff_tail;
wire [0:63] sb_1__0__6_chanx_left_out;
wire [0:63] sb_1__0__6_chanx_right_out;
wire [0:63] sb_1__0__6_chany_top_out;
wire [0:0] sb_1__0__7_ccff_tail;
wire [0:63] sb_1__0__7_chanx_left_out;
wire [0:63] sb_1__0__7_chanx_right_out;
wire [0:63] sb_1__0__7_chany_top_out;
wire [0:0] sb_1__0__8_ccff_tail;
wire [0:63] sb_1__0__8_chanx_left_out;
wire [0:63] sb_1__0__8_chanx_right_out;
wire [0:63] sb_1__0__8_chany_top_out;
wire [0:0] sb_1__18__0_ccff_tail;
wire [0:63] sb_1__18__0_chanx_left_out;
wire [0:63] sb_1__18__0_chanx_right_out;
wire [0:63] sb_1__18__0_chany_bottom_out;
wire [0:0] sb_1__18__1_ccff_tail;
wire [0:63] sb_1__18__1_chanx_left_out;
wire [0:63] sb_1__18__1_chanx_right_out;
wire [0:63] sb_1__18__1_chany_bottom_out;
wire [0:0] sb_1__18__2_ccff_tail;
wire [0:63] sb_1__18__2_chanx_left_out;
wire [0:63] sb_1__18__2_chanx_right_out;
wire [0:63] sb_1__18__2_chany_bottom_out;
wire [0:0] sb_1__18__3_ccff_tail;
wire [0:63] sb_1__18__3_chanx_left_out;
wire [0:63] sb_1__18__3_chanx_right_out;
wire [0:63] sb_1__18__3_chany_bottom_out;
wire [0:0] sb_1__18__4_ccff_tail;
wire [0:63] sb_1__18__4_chanx_left_out;
wire [0:63] sb_1__18__4_chanx_right_out;
wire [0:63] sb_1__18__4_chany_bottom_out;
wire [0:0] sb_1__18__5_ccff_tail;
wire [0:63] sb_1__18__5_chanx_left_out;
wire [0:63] sb_1__18__5_chanx_right_out;
wire [0:63] sb_1__18__5_chany_bottom_out;
wire [0:0] sb_1__18__6_ccff_tail;
wire [0:63] sb_1__18__6_chanx_left_out;
wire [0:63] sb_1__18__6_chanx_right_out;
wire [0:63] sb_1__18__6_chany_bottom_out;
wire [0:0] sb_1__18__7_ccff_tail;
wire [0:63] sb_1__18__7_chanx_left_out;
wire [0:63] sb_1__18__7_chanx_right_out;
wire [0:63] sb_1__18__7_chany_bottom_out;
wire [0:0] sb_1__18__8_ccff_tail;
wire [0:63] sb_1__18__8_chanx_left_out;
wire [0:63] sb_1__18__8_chanx_right_out;
wire [0:63] sb_1__18__8_chany_bottom_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:63] sb_1__1__0_chanx_left_out;
wire [0:63] sb_1__1__0_chanx_right_out;
wire [0:63] sb_1__1__0_chany_bottom_out;
wire [0:63] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__100_ccff_tail;
wire [0:63] sb_1__1__100_chanx_left_out;
wire [0:63] sb_1__1__100_chanx_right_out;
wire [0:63] sb_1__1__100_chany_bottom_out;
wire [0:63] sb_1__1__100_chany_top_out;
wire [0:0] sb_1__1__101_ccff_tail;
wire [0:63] sb_1__1__101_chanx_left_out;
wire [0:63] sb_1__1__101_chanx_right_out;
wire [0:63] sb_1__1__101_chany_bottom_out;
wire [0:63] sb_1__1__101_chany_top_out;
wire [0:0] sb_1__1__102_ccff_tail;
wire [0:63] sb_1__1__102_chanx_left_out;
wire [0:63] sb_1__1__102_chanx_right_out;
wire [0:63] sb_1__1__102_chany_bottom_out;
wire [0:63] sb_1__1__102_chany_top_out;
wire [0:0] sb_1__1__103_ccff_tail;
wire [0:63] sb_1__1__103_chanx_left_out;
wire [0:63] sb_1__1__103_chanx_right_out;
wire [0:63] sb_1__1__103_chany_bottom_out;
wire [0:63] sb_1__1__103_chany_top_out;
wire [0:0] sb_1__1__104_ccff_tail;
wire [0:63] sb_1__1__104_chanx_left_out;
wire [0:63] sb_1__1__104_chanx_right_out;
wire [0:63] sb_1__1__104_chany_bottom_out;
wire [0:63] sb_1__1__104_chany_top_out;
wire [0:0] sb_1__1__105_ccff_tail;
wire [0:63] sb_1__1__105_chanx_left_out;
wire [0:63] sb_1__1__105_chanx_right_out;
wire [0:63] sb_1__1__105_chany_bottom_out;
wire [0:63] sb_1__1__105_chany_top_out;
wire [0:0] sb_1__1__106_ccff_tail;
wire [0:63] sb_1__1__106_chanx_left_out;
wire [0:63] sb_1__1__106_chanx_right_out;
wire [0:63] sb_1__1__106_chany_bottom_out;
wire [0:63] sb_1__1__106_chany_top_out;
wire [0:0] sb_1__1__107_ccff_tail;
wire [0:63] sb_1__1__107_chanx_left_out;
wire [0:63] sb_1__1__107_chanx_right_out;
wire [0:63] sb_1__1__107_chany_bottom_out;
wire [0:63] sb_1__1__107_chany_top_out;
wire [0:0] sb_1__1__108_ccff_tail;
wire [0:63] sb_1__1__108_chanx_left_out;
wire [0:63] sb_1__1__108_chanx_right_out;
wire [0:63] sb_1__1__108_chany_bottom_out;
wire [0:63] sb_1__1__108_chany_top_out;
wire [0:0] sb_1__1__109_ccff_tail;
wire [0:63] sb_1__1__109_chanx_left_out;
wire [0:63] sb_1__1__109_chanx_right_out;
wire [0:63] sb_1__1__109_chany_bottom_out;
wire [0:63] sb_1__1__109_chany_top_out;
wire [0:0] sb_1__1__10_ccff_tail;
wire [0:63] sb_1__1__10_chanx_left_out;
wire [0:63] sb_1__1__10_chanx_right_out;
wire [0:63] sb_1__1__10_chany_bottom_out;
wire [0:63] sb_1__1__10_chany_top_out;
wire [0:0] sb_1__1__110_ccff_tail;
wire [0:63] sb_1__1__110_chanx_left_out;
wire [0:63] sb_1__1__110_chanx_right_out;
wire [0:63] sb_1__1__110_chany_bottom_out;
wire [0:63] sb_1__1__110_chany_top_out;
wire [0:0] sb_1__1__111_ccff_tail;
wire [0:63] sb_1__1__111_chanx_left_out;
wire [0:63] sb_1__1__111_chanx_right_out;
wire [0:63] sb_1__1__111_chany_bottom_out;
wire [0:63] sb_1__1__111_chany_top_out;
wire [0:0] sb_1__1__112_ccff_tail;
wire [0:63] sb_1__1__112_chanx_left_out;
wire [0:63] sb_1__1__112_chanx_right_out;
wire [0:63] sb_1__1__112_chany_bottom_out;
wire [0:63] sb_1__1__112_chany_top_out;
wire [0:0] sb_1__1__113_ccff_tail;
wire [0:63] sb_1__1__113_chanx_left_out;
wire [0:63] sb_1__1__113_chanx_right_out;
wire [0:63] sb_1__1__113_chany_bottom_out;
wire [0:63] sb_1__1__113_chany_top_out;
wire [0:0] sb_1__1__114_ccff_tail;
wire [0:63] sb_1__1__114_chanx_left_out;
wire [0:63] sb_1__1__114_chanx_right_out;
wire [0:63] sb_1__1__114_chany_bottom_out;
wire [0:63] sb_1__1__114_chany_top_out;
wire [0:0] sb_1__1__115_ccff_tail;
wire [0:63] sb_1__1__115_chanx_left_out;
wire [0:63] sb_1__1__115_chanx_right_out;
wire [0:63] sb_1__1__115_chany_bottom_out;
wire [0:63] sb_1__1__115_chany_top_out;
wire [0:0] sb_1__1__116_ccff_tail;
wire [0:63] sb_1__1__116_chanx_left_out;
wire [0:63] sb_1__1__116_chanx_right_out;
wire [0:63] sb_1__1__116_chany_bottom_out;
wire [0:63] sb_1__1__116_chany_top_out;
wire [0:0] sb_1__1__117_ccff_tail;
wire [0:63] sb_1__1__117_chanx_left_out;
wire [0:63] sb_1__1__117_chanx_right_out;
wire [0:63] sb_1__1__117_chany_bottom_out;
wire [0:63] sb_1__1__117_chany_top_out;
wire [0:0] sb_1__1__118_ccff_tail;
wire [0:63] sb_1__1__118_chanx_left_out;
wire [0:63] sb_1__1__118_chanx_right_out;
wire [0:63] sb_1__1__118_chany_bottom_out;
wire [0:63] sb_1__1__118_chany_top_out;
wire [0:0] sb_1__1__119_ccff_tail;
wire [0:63] sb_1__1__119_chanx_left_out;
wire [0:63] sb_1__1__119_chanx_right_out;
wire [0:63] sb_1__1__119_chany_bottom_out;
wire [0:63] sb_1__1__119_chany_top_out;
wire [0:0] sb_1__1__11_ccff_tail;
wire [0:63] sb_1__1__11_chanx_left_out;
wire [0:63] sb_1__1__11_chanx_right_out;
wire [0:63] sb_1__1__11_chany_bottom_out;
wire [0:63] sb_1__1__11_chany_top_out;
wire [0:0] sb_1__1__120_ccff_tail;
wire [0:63] sb_1__1__120_chanx_left_out;
wire [0:63] sb_1__1__120_chanx_right_out;
wire [0:63] sb_1__1__120_chany_bottom_out;
wire [0:63] sb_1__1__120_chany_top_out;
wire [0:0] sb_1__1__121_ccff_tail;
wire [0:63] sb_1__1__121_chanx_left_out;
wire [0:63] sb_1__1__121_chanx_right_out;
wire [0:63] sb_1__1__121_chany_bottom_out;
wire [0:63] sb_1__1__121_chany_top_out;
wire [0:0] sb_1__1__122_ccff_tail;
wire [0:63] sb_1__1__122_chanx_left_out;
wire [0:63] sb_1__1__122_chanx_right_out;
wire [0:63] sb_1__1__122_chany_bottom_out;
wire [0:63] sb_1__1__122_chany_top_out;
wire [0:0] sb_1__1__123_ccff_tail;
wire [0:63] sb_1__1__123_chanx_left_out;
wire [0:63] sb_1__1__123_chanx_right_out;
wire [0:63] sb_1__1__123_chany_bottom_out;
wire [0:63] sb_1__1__123_chany_top_out;
wire [0:0] sb_1__1__124_ccff_tail;
wire [0:63] sb_1__1__124_chanx_left_out;
wire [0:63] sb_1__1__124_chanx_right_out;
wire [0:63] sb_1__1__124_chany_bottom_out;
wire [0:63] sb_1__1__124_chany_top_out;
wire [0:0] sb_1__1__125_ccff_tail;
wire [0:63] sb_1__1__125_chanx_left_out;
wire [0:63] sb_1__1__125_chanx_right_out;
wire [0:63] sb_1__1__125_chany_bottom_out;
wire [0:63] sb_1__1__125_chany_top_out;
wire [0:0] sb_1__1__126_ccff_tail;
wire [0:63] sb_1__1__126_chanx_left_out;
wire [0:63] sb_1__1__126_chanx_right_out;
wire [0:63] sb_1__1__126_chany_bottom_out;
wire [0:63] sb_1__1__126_chany_top_out;
wire [0:0] sb_1__1__127_ccff_tail;
wire [0:63] sb_1__1__127_chanx_left_out;
wire [0:63] sb_1__1__127_chanx_right_out;
wire [0:63] sb_1__1__127_chany_bottom_out;
wire [0:63] sb_1__1__127_chany_top_out;
wire [0:0] sb_1__1__128_ccff_tail;
wire [0:63] sb_1__1__128_chanx_left_out;
wire [0:63] sb_1__1__128_chanx_right_out;
wire [0:63] sb_1__1__128_chany_bottom_out;
wire [0:63] sb_1__1__128_chany_top_out;
wire [0:0] sb_1__1__129_ccff_tail;
wire [0:63] sb_1__1__129_chanx_left_out;
wire [0:63] sb_1__1__129_chanx_right_out;
wire [0:63] sb_1__1__129_chany_bottom_out;
wire [0:63] sb_1__1__129_chany_top_out;
wire [0:0] sb_1__1__12_ccff_tail;
wire [0:63] sb_1__1__12_chanx_left_out;
wire [0:63] sb_1__1__12_chanx_right_out;
wire [0:63] sb_1__1__12_chany_bottom_out;
wire [0:63] sb_1__1__12_chany_top_out;
wire [0:0] sb_1__1__130_ccff_tail;
wire [0:63] sb_1__1__130_chanx_left_out;
wire [0:63] sb_1__1__130_chanx_right_out;
wire [0:63] sb_1__1__130_chany_bottom_out;
wire [0:63] sb_1__1__130_chany_top_out;
wire [0:0] sb_1__1__131_ccff_tail;
wire [0:63] sb_1__1__131_chanx_left_out;
wire [0:63] sb_1__1__131_chanx_right_out;
wire [0:63] sb_1__1__131_chany_bottom_out;
wire [0:63] sb_1__1__131_chany_top_out;
wire [0:0] sb_1__1__132_ccff_tail;
wire [0:63] sb_1__1__132_chanx_left_out;
wire [0:63] sb_1__1__132_chanx_right_out;
wire [0:63] sb_1__1__132_chany_bottom_out;
wire [0:63] sb_1__1__132_chany_top_out;
wire [0:0] sb_1__1__133_ccff_tail;
wire [0:63] sb_1__1__133_chanx_left_out;
wire [0:63] sb_1__1__133_chanx_right_out;
wire [0:63] sb_1__1__133_chany_bottom_out;
wire [0:63] sb_1__1__133_chany_top_out;
wire [0:0] sb_1__1__134_ccff_tail;
wire [0:63] sb_1__1__134_chanx_left_out;
wire [0:63] sb_1__1__134_chanx_right_out;
wire [0:63] sb_1__1__134_chany_bottom_out;
wire [0:63] sb_1__1__134_chany_top_out;
wire [0:0] sb_1__1__135_ccff_tail;
wire [0:63] sb_1__1__135_chanx_left_out;
wire [0:63] sb_1__1__135_chanx_right_out;
wire [0:63] sb_1__1__135_chany_bottom_out;
wire [0:63] sb_1__1__135_chany_top_out;
wire [0:0] sb_1__1__136_ccff_tail;
wire [0:63] sb_1__1__136_chanx_left_out;
wire [0:63] sb_1__1__136_chanx_right_out;
wire [0:63] sb_1__1__136_chany_bottom_out;
wire [0:63] sb_1__1__136_chany_top_out;
wire [0:0] sb_1__1__137_ccff_tail;
wire [0:63] sb_1__1__137_chanx_left_out;
wire [0:63] sb_1__1__137_chanx_right_out;
wire [0:63] sb_1__1__137_chany_bottom_out;
wire [0:63] sb_1__1__137_chany_top_out;
wire [0:0] sb_1__1__138_ccff_tail;
wire [0:63] sb_1__1__138_chanx_left_out;
wire [0:63] sb_1__1__138_chanx_right_out;
wire [0:63] sb_1__1__138_chany_bottom_out;
wire [0:63] sb_1__1__138_chany_top_out;
wire [0:0] sb_1__1__139_ccff_tail;
wire [0:63] sb_1__1__139_chanx_left_out;
wire [0:63] sb_1__1__139_chanx_right_out;
wire [0:63] sb_1__1__139_chany_bottom_out;
wire [0:63] sb_1__1__139_chany_top_out;
wire [0:0] sb_1__1__13_ccff_tail;
wire [0:63] sb_1__1__13_chanx_left_out;
wire [0:63] sb_1__1__13_chanx_right_out;
wire [0:63] sb_1__1__13_chany_bottom_out;
wire [0:63] sb_1__1__13_chany_top_out;
wire [0:0] sb_1__1__140_ccff_tail;
wire [0:63] sb_1__1__140_chanx_left_out;
wire [0:63] sb_1__1__140_chanx_right_out;
wire [0:63] sb_1__1__140_chany_bottom_out;
wire [0:63] sb_1__1__140_chany_top_out;
wire [0:0] sb_1__1__141_ccff_tail;
wire [0:63] sb_1__1__141_chanx_left_out;
wire [0:63] sb_1__1__141_chanx_right_out;
wire [0:63] sb_1__1__141_chany_bottom_out;
wire [0:63] sb_1__1__141_chany_top_out;
wire [0:0] sb_1__1__142_ccff_tail;
wire [0:63] sb_1__1__142_chanx_left_out;
wire [0:63] sb_1__1__142_chanx_right_out;
wire [0:63] sb_1__1__142_chany_bottom_out;
wire [0:63] sb_1__1__142_chany_top_out;
wire [0:0] sb_1__1__143_ccff_tail;
wire [0:63] sb_1__1__143_chanx_left_out;
wire [0:63] sb_1__1__143_chanx_right_out;
wire [0:63] sb_1__1__143_chany_bottom_out;
wire [0:63] sb_1__1__143_chany_top_out;
wire [0:0] sb_1__1__144_ccff_tail;
wire [0:63] sb_1__1__144_chanx_left_out;
wire [0:63] sb_1__1__144_chanx_right_out;
wire [0:63] sb_1__1__144_chany_bottom_out;
wire [0:63] sb_1__1__144_chany_top_out;
wire [0:0] sb_1__1__145_ccff_tail;
wire [0:63] sb_1__1__145_chanx_left_out;
wire [0:63] sb_1__1__145_chanx_right_out;
wire [0:63] sb_1__1__145_chany_bottom_out;
wire [0:63] sb_1__1__145_chany_top_out;
wire [0:63] sb_1__1__146_chanx_left_out;
wire [0:63] sb_1__1__146_chanx_right_out;
wire [0:63] sb_1__1__146_chany_bottom_out;
wire [0:63] sb_1__1__146_chany_top_out;
wire [0:0] sb_1__1__147_ccff_tail;
wire [0:63] sb_1__1__147_chanx_left_out;
wire [0:63] sb_1__1__147_chanx_right_out;
wire [0:63] sb_1__1__147_chany_bottom_out;
wire [0:63] sb_1__1__147_chany_top_out;
wire [0:0] sb_1__1__148_ccff_tail;
wire [0:63] sb_1__1__148_chanx_left_out;
wire [0:63] sb_1__1__148_chanx_right_out;
wire [0:63] sb_1__1__148_chany_bottom_out;
wire [0:63] sb_1__1__148_chany_top_out;
wire [0:0] sb_1__1__149_ccff_tail;
wire [0:63] sb_1__1__149_chanx_left_out;
wire [0:63] sb_1__1__149_chanx_right_out;
wire [0:63] sb_1__1__149_chany_bottom_out;
wire [0:63] sb_1__1__149_chany_top_out;
wire [0:0] sb_1__1__14_ccff_tail;
wire [0:63] sb_1__1__14_chanx_left_out;
wire [0:63] sb_1__1__14_chanx_right_out;
wire [0:63] sb_1__1__14_chany_bottom_out;
wire [0:63] sb_1__1__14_chany_top_out;
wire [0:0] sb_1__1__150_ccff_tail;
wire [0:63] sb_1__1__150_chanx_left_out;
wire [0:63] sb_1__1__150_chanx_right_out;
wire [0:63] sb_1__1__150_chany_bottom_out;
wire [0:63] sb_1__1__150_chany_top_out;
wire [0:0] sb_1__1__151_ccff_tail;
wire [0:63] sb_1__1__151_chanx_left_out;
wire [0:63] sb_1__1__151_chanx_right_out;
wire [0:63] sb_1__1__151_chany_bottom_out;
wire [0:63] sb_1__1__151_chany_top_out;
wire [0:0] sb_1__1__152_ccff_tail;
wire [0:63] sb_1__1__152_chanx_left_out;
wire [0:63] sb_1__1__152_chanx_right_out;
wire [0:63] sb_1__1__152_chany_bottom_out;
wire [0:63] sb_1__1__152_chany_top_out;
wire [0:0] sb_1__1__15_ccff_tail;
wire [0:63] sb_1__1__15_chanx_left_out;
wire [0:63] sb_1__1__15_chanx_right_out;
wire [0:63] sb_1__1__15_chany_bottom_out;
wire [0:63] sb_1__1__15_chany_top_out;
wire [0:0] sb_1__1__16_ccff_tail;
wire [0:63] sb_1__1__16_chanx_left_out;
wire [0:63] sb_1__1__16_chanx_right_out;
wire [0:63] sb_1__1__16_chany_bottom_out;
wire [0:63] sb_1__1__16_chany_top_out;
wire [0:0] sb_1__1__17_ccff_tail;
wire [0:63] sb_1__1__17_chanx_left_out;
wire [0:63] sb_1__1__17_chanx_right_out;
wire [0:63] sb_1__1__17_chany_bottom_out;
wire [0:63] sb_1__1__17_chany_top_out;
wire [0:0] sb_1__1__18_ccff_tail;
wire [0:63] sb_1__1__18_chanx_left_out;
wire [0:63] sb_1__1__18_chanx_right_out;
wire [0:63] sb_1__1__18_chany_bottom_out;
wire [0:63] sb_1__1__18_chany_top_out;
wire [0:0] sb_1__1__19_ccff_tail;
wire [0:63] sb_1__1__19_chanx_left_out;
wire [0:63] sb_1__1__19_chanx_right_out;
wire [0:63] sb_1__1__19_chany_bottom_out;
wire [0:63] sb_1__1__19_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:63] sb_1__1__1_chanx_left_out;
wire [0:63] sb_1__1__1_chanx_right_out;
wire [0:63] sb_1__1__1_chany_bottom_out;
wire [0:63] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__20_ccff_tail;
wire [0:63] sb_1__1__20_chanx_left_out;
wire [0:63] sb_1__1__20_chanx_right_out;
wire [0:63] sb_1__1__20_chany_bottom_out;
wire [0:63] sb_1__1__20_chany_top_out;
wire [0:0] sb_1__1__21_ccff_tail;
wire [0:63] sb_1__1__21_chanx_left_out;
wire [0:63] sb_1__1__21_chanx_right_out;
wire [0:63] sb_1__1__21_chany_bottom_out;
wire [0:63] sb_1__1__21_chany_top_out;
wire [0:0] sb_1__1__22_ccff_tail;
wire [0:63] sb_1__1__22_chanx_left_out;
wire [0:63] sb_1__1__22_chanx_right_out;
wire [0:63] sb_1__1__22_chany_bottom_out;
wire [0:63] sb_1__1__22_chany_top_out;
wire [0:0] sb_1__1__23_ccff_tail;
wire [0:63] sb_1__1__23_chanx_left_out;
wire [0:63] sb_1__1__23_chanx_right_out;
wire [0:63] sb_1__1__23_chany_bottom_out;
wire [0:63] sb_1__1__23_chany_top_out;
wire [0:0] sb_1__1__24_ccff_tail;
wire [0:63] sb_1__1__24_chanx_left_out;
wire [0:63] sb_1__1__24_chanx_right_out;
wire [0:63] sb_1__1__24_chany_bottom_out;
wire [0:63] sb_1__1__24_chany_top_out;
wire [0:0] sb_1__1__25_ccff_tail;
wire [0:63] sb_1__1__25_chanx_left_out;
wire [0:63] sb_1__1__25_chanx_right_out;
wire [0:63] sb_1__1__25_chany_bottom_out;
wire [0:63] sb_1__1__25_chany_top_out;
wire [0:0] sb_1__1__26_ccff_tail;
wire [0:63] sb_1__1__26_chanx_left_out;
wire [0:63] sb_1__1__26_chanx_right_out;
wire [0:63] sb_1__1__26_chany_bottom_out;
wire [0:63] sb_1__1__26_chany_top_out;
wire [0:0] sb_1__1__27_ccff_tail;
wire [0:63] sb_1__1__27_chanx_left_out;
wire [0:63] sb_1__1__27_chanx_right_out;
wire [0:63] sb_1__1__27_chany_bottom_out;
wire [0:63] sb_1__1__27_chany_top_out;
wire [0:0] sb_1__1__28_ccff_tail;
wire [0:63] sb_1__1__28_chanx_left_out;
wire [0:63] sb_1__1__28_chanx_right_out;
wire [0:63] sb_1__1__28_chany_bottom_out;
wire [0:63] sb_1__1__28_chany_top_out;
wire [0:0] sb_1__1__29_ccff_tail;
wire [0:63] sb_1__1__29_chanx_left_out;
wire [0:63] sb_1__1__29_chanx_right_out;
wire [0:63] sb_1__1__29_chany_bottom_out;
wire [0:63] sb_1__1__29_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:63] sb_1__1__2_chanx_left_out;
wire [0:63] sb_1__1__2_chanx_right_out;
wire [0:63] sb_1__1__2_chany_bottom_out;
wire [0:63] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__30_ccff_tail;
wire [0:63] sb_1__1__30_chanx_left_out;
wire [0:63] sb_1__1__30_chanx_right_out;
wire [0:63] sb_1__1__30_chany_bottom_out;
wire [0:63] sb_1__1__30_chany_top_out;
wire [0:0] sb_1__1__31_ccff_tail;
wire [0:63] sb_1__1__31_chanx_left_out;
wire [0:63] sb_1__1__31_chanx_right_out;
wire [0:63] sb_1__1__31_chany_bottom_out;
wire [0:63] sb_1__1__31_chany_top_out;
wire [0:0] sb_1__1__32_ccff_tail;
wire [0:63] sb_1__1__32_chanx_left_out;
wire [0:63] sb_1__1__32_chanx_right_out;
wire [0:63] sb_1__1__32_chany_bottom_out;
wire [0:63] sb_1__1__32_chany_top_out;
wire [0:0] sb_1__1__33_ccff_tail;
wire [0:63] sb_1__1__33_chanx_left_out;
wire [0:63] sb_1__1__33_chanx_right_out;
wire [0:63] sb_1__1__33_chany_bottom_out;
wire [0:63] sb_1__1__33_chany_top_out;
wire [0:0] sb_1__1__34_ccff_tail;
wire [0:63] sb_1__1__34_chanx_left_out;
wire [0:63] sb_1__1__34_chanx_right_out;
wire [0:63] sb_1__1__34_chany_bottom_out;
wire [0:63] sb_1__1__34_chany_top_out;
wire [0:0] sb_1__1__35_ccff_tail;
wire [0:63] sb_1__1__35_chanx_left_out;
wire [0:63] sb_1__1__35_chanx_right_out;
wire [0:63] sb_1__1__35_chany_bottom_out;
wire [0:63] sb_1__1__35_chany_top_out;
wire [0:0] sb_1__1__36_ccff_tail;
wire [0:63] sb_1__1__36_chanx_left_out;
wire [0:63] sb_1__1__36_chanx_right_out;
wire [0:63] sb_1__1__36_chany_bottom_out;
wire [0:63] sb_1__1__36_chany_top_out;
wire [0:0] sb_1__1__37_ccff_tail;
wire [0:63] sb_1__1__37_chanx_left_out;
wire [0:63] sb_1__1__37_chanx_right_out;
wire [0:63] sb_1__1__37_chany_bottom_out;
wire [0:63] sb_1__1__37_chany_top_out;
wire [0:0] sb_1__1__38_ccff_tail;
wire [0:63] sb_1__1__38_chanx_left_out;
wire [0:63] sb_1__1__38_chanx_right_out;
wire [0:63] sb_1__1__38_chany_bottom_out;
wire [0:63] sb_1__1__38_chany_top_out;
wire [0:0] sb_1__1__39_ccff_tail;
wire [0:63] sb_1__1__39_chanx_left_out;
wire [0:63] sb_1__1__39_chanx_right_out;
wire [0:63] sb_1__1__39_chany_bottom_out;
wire [0:63] sb_1__1__39_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:63] sb_1__1__3_chanx_left_out;
wire [0:63] sb_1__1__3_chanx_right_out;
wire [0:63] sb_1__1__3_chany_bottom_out;
wire [0:63] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__40_ccff_tail;
wire [0:63] sb_1__1__40_chanx_left_out;
wire [0:63] sb_1__1__40_chanx_right_out;
wire [0:63] sb_1__1__40_chany_bottom_out;
wire [0:63] sb_1__1__40_chany_top_out;
wire [0:0] sb_1__1__41_ccff_tail;
wire [0:63] sb_1__1__41_chanx_left_out;
wire [0:63] sb_1__1__41_chanx_right_out;
wire [0:63] sb_1__1__41_chany_bottom_out;
wire [0:63] sb_1__1__41_chany_top_out;
wire [0:0] sb_1__1__42_ccff_tail;
wire [0:63] sb_1__1__42_chanx_left_out;
wire [0:63] sb_1__1__42_chanx_right_out;
wire [0:63] sb_1__1__42_chany_bottom_out;
wire [0:63] sb_1__1__42_chany_top_out;
wire [0:0] sb_1__1__43_ccff_tail;
wire [0:63] sb_1__1__43_chanx_left_out;
wire [0:63] sb_1__1__43_chanx_right_out;
wire [0:63] sb_1__1__43_chany_bottom_out;
wire [0:63] sb_1__1__43_chany_top_out;
wire [0:0] sb_1__1__44_ccff_tail;
wire [0:63] sb_1__1__44_chanx_left_out;
wire [0:63] sb_1__1__44_chanx_right_out;
wire [0:63] sb_1__1__44_chany_bottom_out;
wire [0:63] sb_1__1__44_chany_top_out;
wire [0:0] sb_1__1__45_ccff_tail;
wire [0:63] sb_1__1__45_chanx_left_out;
wire [0:63] sb_1__1__45_chanx_right_out;
wire [0:63] sb_1__1__45_chany_bottom_out;
wire [0:63] sb_1__1__45_chany_top_out;
wire [0:0] sb_1__1__46_ccff_tail;
wire [0:63] sb_1__1__46_chanx_left_out;
wire [0:63] sb_1__1__46_chanx_right_out;
wire [0:63] sb_1__1__46_chany_bottom_out;
wire [0:63] sb_1__1__46_chany_top_out;
wire [0:0] sb_1__1__47_ccff_tail;
wire [0:63] sb_1__1__47_chanx_left_out;
wire [0:63] sb_1__1__47_chanx_right_out;
wire [0:63] sb_1__1__47_chany_bottom_out;
wire [0:63] sb_1__1__47_chany_top_out;
wire [0:0] sb_1__1__48_ccff_tail;
wire [0:63] sb_1__1__48_chanx_left_out;
wire [0:63] sb_1__1__48_chanx_right_out;
wire [0:63] sb_1__1__48_chany_bottom_out;
wire [0:63] sb_1__1__48_chany_top_out;
wire [0:0] sb_1__1__49_ccff_tail;
wire [0:63] sb_1__1__49_chanx_left_out;
wire [0:63] sb_1__1__49_chanx_right_out;
wire [0:63] sb_1__1__49_chany_bottom_out;
wire [0:63] sb_1__1__49_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:63] sb_1__1__4_chanx_left_out;
wire [0:63] sb_1__1__4_chanx_right_out;
wire [0:63] sb_1__1__4_chany_bottom_out;
wire [0:63] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__50_ccff_tail;
wire [0:63] sb_1__1__50_chanx_left_out;
wire [0:63] sb_1__1__50_chanx_right_out;
wire [0:63] sb_1__1__50_chany_bottom_out;
wire [0:63] sb_1__1__50_chany_top_out;
wire [0:0] sb_1__1__51_ccff_tail;
wire [0:63] sb_1__1__51_chanx_left_out;
wire [0:63] sb_1__1__51_chanx_right_out;
wire [0:63] sb_1__1__51_chany_bottom_out;
wire [0:63] sb_1__1__51_chany_top_out;
wire [0:0] sb_1__1__52_ccff_tail;
wire [0:63] sb_1__1__52_chanx_left_out;
wire [0:63] sb_1__1__52_chanx_right_out;
wire [0:63] sb_1__1__52_chany_bottom_out;
wire [0:63] sb_1__1__52_chany_top_out;
wire [0:0] sb_1__1__53_ccff_tail;
wire [0:63] sb_1__1__53_chanx_left_out;
wire [0:63] sb_1__1__53_chanx_right_out;
wire [0:63] sb_1__1__53_chany_bottom_out;
wire [0:63] sb_1__1__53_chany_top_out;
wire [0:0] sb_1__1__54_ccff_tail;
wire [0:63] sb_1__1__54_chanx_left_out;
wire [0:63] sb_1__1__54_chanx_right_out;
wire [0:63] sb_1__1__54_chany_bottom_out;
wire [0:63] sb_1__1__54_chany_top_out;
wire [0:0] sb_1__1__55_ccff_tail;
wire [0:63] sb_1__1__55_chanx_left_out;
wire [0:63] sb_1__1__55_chanx_right_out;
wire [0:63] sb_1__1__55_chany_bottom_out;
wire [0:63] sb_1__1__55_chany_top_out;
wire [0:0] sb_1__1__56_ccff_tail;
wire [0:63] sb_1__1__56_chanx_left_out;
wire [0:63] sb_1__1__56_chanx_right_out;
wire [0:63] sb_1__1__56_chany_bottom_out;
wire [0:63] sb_1__1__56_chany_top_out;
wire [0:0] sb_1__1__57_ccff_tail;
wire [0:63] sb_1__1__57_chanx_left_out;
wire [0:63] sb_1__1__57_chanx_right_out;
wire [0:63] sb_1__1__57_chany_bottom_out;
wire [0:63] sb_1__1__57_chany_top_out;
wire [0:0] sb_1__1__58_ccff_tail;
wire [0:63] sb_1__1__58_chanx_left_out;
wire [0:63] sb_1__1__58_chanx_right_out;
wire [0:63] sb_1__1__58_chany_bottom_out;
wire [0:63] sb_1__1__58_chany_top_out;
wire [0:0] sb_1__1__59_ccff_tail;
wire [0:63] sb_1__1__59_chanx_left_out;
wire [0:63] sb_1__1__59_chanx_right_out;
wire [0:63] sb_1__1__59_chany_bottom_out;
wire [0:63] sb_1__1__59_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:63] sb_1__1__5_chanx_left_out;
wire [0:63] sb_1__1__5_chanx_right_out;
wire [0:63] sb_1__1__5_chany_bottom_out;
wire [0:63] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__60_ccff_tail;
wire [0:63] sb_1__1__60_chanx_left_out;
wire [0:63] sb_1__1__60_chanx_right_out;
wire [0:63] sb_1__1__60_chany_bottom_out;
wire [0:63] sb_1__1__60_chany_top_out;
wire [0:0] sb_1__1__61_ccff_tail;
wire [0:63] sb_1__1__61_chanx_left_out;
wire [0:63] sb_1__1__61_chanx_right_out;
wire [0:63] sb_1__1__61_chany_bottom_out;
wire [0:63] sb_1__1__61_chany_top_out;
wire [0:0] sb_1__1__62_ccff_tail;
wire [0:63] sb_1__1__62_chanx_left_out;
wire [0:63] sb_1__1__62_chanx_right_out;
wire [0:63] sb_1__1__62_chany_bottom_out;
wire [0:63] sb_1__1__62_chany_top_out;
wire [0:0] sb_1__1__63_ccff_tail;
wire [0:63] sb_1__1__63_chanx_left_out;
wire [0:63] sb_1__1__63_chanx_right_out;
wire [0:63] sb_1__1__63_chany_bottom_out;
wire [0:63] sb_1__1__63_chany_top_out;
wire [0:0] sb_1__1__64_ccff_tail;
wire [0:63] sb_1__1__64_chanx_left_out;
wire [0:63] sb_1__1__64_chanx_right_out;
wire [0:63] sb_1__1__64_chany_bottom_out;
wire [0:63] sb_1__1__64_chany_top_out;
wire [0:0] sb_1__1__65_ccff_tail;
wire [0:63] sb_1__1__65_chanx_left_out;
wire [0:63] sb_1__1__65_chanx_right_out;
wire [0:63] sb_1__1__65_chany_bottom_out;
wire [0:63] sb_1__1__65_chany_top_out;
wire [0:0] sb_1__1__66_ccff_tail;
wire [0:63] sb_1__1__66_chanx_left_out;
wire [0:63] sb_1__1__66_chanx_right_out;
wire [0:63] sb_1__1__66_chany_bottom_out;
wire [0:63] sb_1__1__66_chany_top_out;
wire [0:0] sb_1__1__67_ccff_tail;
wire [0:63] sb_1__1__67_chanx_left_out;
wire [0:63] sb_1__1__67_chanx_right_out;
wire [0:63] sb_1__1__67_chany_bottom_out;
wire [0:63] sb_1__1__67_chany_top_out;
wire [0:0] sb_1__1__68_ccff_tail;
wire [0:63] sb_1__1__68_chanx_left_out;
wire [0:63] sb_1__1__68_chanx_right_out;
wire [0:63] sb_1__1__68_chany_bottom_out;
wire [0:63] sb_1__1__68_chany_top_out;
wire [0:0] sb_1__1__69_ccff_tail;
wire [0:63] sb_1__1__69_chanx_left_out;
wire [0:63] sb_1__1__69_chanx_right_out;
wire [0:63] sb_1__1__69_chany_bottom_out;
wire [0:63] sb_1__1__69_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:63] sb_1__1__6_chanx_left_out;
wire [0:63] sb_1__1__6_chanx_right_out;
wire [0:63] sb_1__1__6_chany_bottom_out;
wire [0:63] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__70_ccff_tail;
wire [0:63] sb_1__1__70_chanx_left_out;
wire [0:63] sb_1__1__70_chanx_right_out;
wire [0:63] sb_1__1__70_chany_bottom_out;
wire [0:63] sb_1__1__70_chany_top_out;
wire [0:0] sb_1__1__71_ccff_tail;
wire [0:63] sb_1__1__71_chanx_left_out;
wire [0:63] sb_1__1__71_chanx_right_out;
wire [0:63] sb_1__1__71_chany_bottom_out;
wire [0:63] sb_1__1__71_chany_top_out;
wire [0:0] sb_1__1__72_ccff_tail;
wire [0:63] sb_1__1__72_chanx_left_out;
wire [0:63] sb_1__1__72_chanx_right_out;
wire [0:63] sb_1__1__72_chany_bottom_out;
wire [0:63] sb_1__1__72_chany_top_out;
wire [0:0] sb_1__1__73_ccff_tail;
wire [0:63] sb_1__1__73_chanx_left_out;
wire [0:63] sb_1__1__73_chanx_right_out;
wire [0:63] sb_1__1__73_chany_bottom_out;
wire [0:63] sb_1__1__73_chany_top_out;
wire [0:0] sb_1__1__74_ccff_tail;
wire [0:63] sb_1__1__74_chanx_left_out;
wire [0:63] sb_1__1__74_chanx_right_out;
wire [0:63] sb_1__1__74_chany_bottom_out;
wire [0:63] sb_1__1__74_chany_top_out;
wire [0:0] sb_1__1__75_ccff_tail;
wire [0:63] sb_1__1__75_chanx_left_out;
wire [0:63] sb_1__1__75_chanx_right_out;
wire [0:63] sb_1__1__75_chany_bottom_out;
wire [0:63] sb_1__1__75_chany_top_out;
wire [0:0] sb_1__1__76_ccff_tail;
wire [0:63] sb_1__1__76_chanx_left_out;
wire [0:63] sb_1__1__76_chanx_right_out;
wire [0:63] sb_1__1__76_chany_bottom_out;
wire [0:63] sb_1__1__76_chany_top_out;
wire [0:0] sb_1__1__77_ccff_tail;
wire [0:63] sb_1__1__77_chanx_left_out;
wire [0:63] sb_1__1__77_chanx_right_out;
wire [0:63] sb_1__1__77_chany_bottom_out;
wire [0:63] sb_1__1__77_chany_top_out;
wire [0:0] sb_1__1__78_ccff_tail;
wire [0:63] sb_1__1__78_chanx_left_out;
wire [0:63] sb_1__1__78_chanx_right_out;
wire [0:63] sb_1__1__78_chany_bottom_out;
wire [0:63] sb_1__1__78_chany_top_out;
wire [0:0] sb_1__1__79_ccff_tail;
wire [0:63] sb_1__1__79_chanx_left_out;
wire [0:63] sb_1__1__79_chanx_right_out;
wire [0:63] sb_1__1__79_chany_bottom_out;
wire [0:63] sb_1__1__79_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:63] sb_1__1__7_chanx_left_out;
wire [0:63] sb_1__1__7_chanx_right_out;
wire [0:63] sb_1__1__7_chany_bottom_out;
wire [0:63] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__80_ccff_tail;
wire [0:63] sb_1__1__80_chanx_left_out;
wire [0:63] sb_1__1__80_chanx_right_out;
wire [0:63] sb_1__1__80_chany_bottom_out;
wire [0:63] sb_1__1__80_chany_top_out;
wire [0:0] sb_1__1__81_ccff_tail;
wire [0:63] sb_1__1__81_chanx_left_out;
wire [0:63] sb_1__1__81_chanx_right_out;
wire [0:63] sb_1__1__81_chany_bottom_out;
wire [0:63] sb_1__1__81_chany_top_out;
wire [0:0] sb_1__1__82_ccff_tail;
wire [0:63] sb_1__1__82_chanx_left_out;
wire [0:63] sb_1__1__82_chanx_right_out;
wire [0:63] sb_1__1__82_chany_bottom_out;
wire [0:63] sb_1__1__82_chany_top_out;
wire [0:0] sb_1__1__83_ccff_tail;
wire [0:63] sb_1__1__83_chanx_left_out;
wire [0:63] sb_1__1__83_chanx_right_out;
wire [0:63] sb_1__1__83_chany_bottom_out;
wire [0:63] sb_1__1__83_chany_top_out;
wire [0:0] sb_1__1__84_ccff_tail;
wire [0:63] sb_1__1__84_chanx_left_out;
wire [0:63] sb_1__1__84_chanx_right_out;
wire [0:63] sb_1__1__84_chany_bottom_out;
wire [0:63] sb_1__1__84_chany_top_out;
wire [0:0] sb_1__1__85_ccff_tail;
wire [0:63] sb_1__1__85_chanx_left_out;
wire [0:63] sb_1__1__85_chanx_right_out;
wire [0:63] sb_1__1__85_chany_bottom_out;
wire [0:63] sb_1__1__85_chany_top_out;
wire [0:0] sb_1__1__86_ccff_tail;
wire [0:63] sb_1__1__86_chanx_left_out;
wire [0:63] sb_1__1__86_chanx_right_out;
wire [0:63] sb_1__1__86_chany_bottom_out;
wire [0:63] sb_1__1__86_chany_top_out;
wire [0:0] sb_1__1__87_ccff_tail;
wire [0:63] sb_1__1__87_chanx_left_out;
wire [0:63] sb_1__1__87_chanx_right_out;
wire [0:63] sb_1__1__87_chany_bottom_out;
wire [0:63] sb_1__1__87_chany_top_out;
wire [0:0] sb_1__1__88_ccff_tail;
wire [0:63] sb_1__1__88_chanx_left_out;
wire [0:63] sb_1__1__88_chanx_right_out;
wire [0:63] sb_1__1__88_chany_bottom_out;
wire [0:63] sb_1__1__88_chany_top_out;
wire [0:0] sb_1__1__89_ccff_tail;
wire [0:63] sb_1__1__89_chanx_left_out;
wire [0:63] sb_1__1__89_chanx_right_out;
wire [0:63] sb_1__1__89_chany_bottom_out;
wire [0:63] sb_1__1__89_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:63] sb_1__1__8_chanx_left_out;
wire [0:63] sb_1__1__8_chanx_right_out;
wire [0:63] sb_1__1__8_chany_bottom_out;
wire [0:63] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__1__90_ccff_tail;
wire [0:63] sb_1__1__90_chanx_left_out;
wire [0:63] sb_1__1__90_chanx_right_out;
wire [0:63] sb_1__1__90_chany_bottom_out;
wire [0:63] sb_1__1__90_chany_top_out;
wire [0:0] sb_1__1__91_ccff_tail;
wire [0:63] sb_1__1__91_chanx_left_out;
wire [0:63] sb_1__1__91_chanx_right_out;
wire [0:63] sb_1__1__91_chany_bottom_out;
wire [0:63] sb_1__1__91_chany_top_out;
wire [0:0] sb_1__1__92_ccff_tail;
wire [0:63] sb_1__1__92_chanx_left_out;
wire [0:63] sb_1__1__92_chanx_right_out;
wire [0:63] sb_1__1__92_chany_bottom_out;
wire [0:63] sb_1__1__92_chany_top_out;
wire [0:0] sb_1__1__93_ccff_tail;
wire [0:63] sb_1__1__93_chanx_left_out;
wire [0:63] sb_1__1__93_chanx_right_out;
wire [0:63] sb_1__1__93_chany_bottom_out;
wire [0:63] sb_1__1__93_chany_top_out;
wire [0:0] sb_1__1__94_ccff_tail;
wire [0:63] sb_1__1__94_chanx_left_out;
wire [0:63] sb_1__1__94_chanx_right_out;
wire [0:63] sb_1__1__94_chany_bottom_out;
wire [0:63] sb_1__1__94_chany_top_out;
wire [0:0] sb_1__1__95_ccff_tail;
wire [0:63] sb_1__1__95_chanx_left_out;
wire [0:63] sb_1__1__95_chanx_right_out;
wire [0:63] sb_1__1__95_chany_bottom_out;
wire [0:63] sb_1__1__95_chany_top_out;
wire [0:0] sb_1__1__96_ccff_tail;
wire [0:63] sb_1__1__96_chanx_left_out;
wire [0:63] sb_1__1__96_chanx_right_out;
wire [0:63] sb_1__1__96_chany_bottom_out;
wire [0:63] sb_1__1__96_chany_top_out;
wire [0:0] sb_1__1__97_ccff_tail;
wire [0:63] sb_1__1__97_chanx_left_out;
wire [0:63] sb_1__1__97_chanx_right_out;
wire [0:63] sb_1__1__97_chany_bottom_out;
wire [0:63] sb_1__1__97_chany_top_out;
wire [0:0] sb_1__1__98_ccff_tail;
wire [0:63] sb_1__1__98_chanx_left_out;
wire [0:63] sb_1__1__98_chanx_right_out;
wire [0:63] sb_1__1__98_chany_bottom_out;
wire [0:63] sb_1__1__98_chany_top_out;
wire [0:0] sb_1__1__99_ccff_tail;
wire [0:63] sb_1__1__99_chanx_left_out;
wire [0:63] sb_1__1__99_chanx_right_out;
wire [0:63] sb_1__1__99_chany_bottom_out;
wire [0:63] sb_1__1__99_chany_top_out;
wire [0:0] sb_1__1__9_ccff_tail;
wire [0:63] sb_1__1__9_chanx_left_out;
wire [0:63] sb_1__1__9_chanx_right_out;
wire [0:63] sb_1__1__9_chany_bottom_out;
wire [0:63] sb_1__1__9_chany_top_out;
wire [0:0] sb_3__0__0_ccff_tail;
wire [0:63] sb_3__0__0_chanx_left_out;
wire [0:63] sb_3__0__0_chanx_right_out;
wire [0:63] sb_3__0__0_chany_top_out;
wire [0:0] sb_3__0__1_ccff_tail;
wire [0:63] sb_3__0__1_chanx_left_out;
wire [0:63] sb_3__0__1_chanx_right_out;
wire [0:63] sb_3__0__1_chany_top_out;
wire [0:0] sb_3__18__0_ccff_tail;
wire [0:63] sb_3__18__0_chanx_left_out;
wire [0:63] sb_3__18__0_chanx_right_out;
wire [0:63] sb_3__18__0_chany_bottom_out;
wire [0:0] sb_3__18__1_ccff_tail;
wire [0:63] sb_3__18__1_chanx_left_out;
wire [0:63] sb_3__18__1_chanx_right_out;
wire [0:63] sb_3__18__1_chany_bottom_out;
wire [0:0] sb_3__1__0_ccff_tail;
wire [0:63] sb_3__1__0_chanx_left_out;
wire [0:63] sb_3__1__0_chanx_right_out;
wire [0:63] sb_3__1__0_chany_bottom_out;
wire [0:63] sb_3__1__0_chany_top_out;
wire [0:0] sb_3__1__10_ccff_tail;
wire [0:63] sb_3__1__10_chanx_left_out;
wire [0:63] sb_3__1__10_chanx_right_out;
wire [0:63] sb_3__1__10_chany_bottom_out;
wire [0:63] sb_3__1__10_chany_top_out;
wire [0:0] sb_3__1__11_ccff_tail;
wire [0:63] sb_3__1__11_chanx_left_out;
wire [0:63] sb_3__1__11_chanx_right_out;
wire [0:63] sb_3__1__11_chany_bottom_out;
wire [0:63] sb_3__1__11_chany_top_out;
wire [0:0] sb_3__1__12_ccff_tail;
wire [0:63] sb_3__1__12_chanx_left_out;
wire [0:63] sb_3__1__12_chanx_right_out;
wire [0:63] sb_3__1__12_chany_bottom_out;
wire [0:63] sb_3__1__12_chany_top_out;
wire [0:0] sb_3__1__13_ccff_tail;
wire [0:63] sb_3__1__13_chanx_left_out;
wire [0:63] sb_3__1__13_chanx_right_out;
wire [0:63] sb_3__1__13_chany_bottom_out;
wire [0:63] sb_3__1__13_chany_top_out;
wire [0:0] sb_3__1__14_ccff_tail;
wire [0:63] sb_3__1__14_chanx_left_out;
wire [0:63] sb_3__1__14_chanx_right_out;
wire [0:63] sb_3__1__14_chany_bottom_out;
wire [0:63] sb_3__1__14_chany_top_out;
wire [0:0] sb_3__1__15_ccff_tail;
wire [0:63] sb_3__1__15_chanx_left_out;
wire [0:63] sb_3__1__15_chanx_right_out;
wire [0:63] sb_3__1__15_chany_bottom_out;
wire [0:63] sb_3__1__15_chany_top_out;
wire [0:0] sb_3__1__16_ccff_tail;
wire [0:63] sb_3__1__16_chanx_left_out;
wire [0:63] sb_3__1__16_chanx_right_out;
wire [0:63] sb_3__1__16_chany_bottom_out;
wire [0:63] sb_3__1__16_chany_top_out;
wire [0:0] sb_3__1__17_ccff_tail;
wire [0:63] sb_3__1__17_chanx_left_out;
wire [0:63] sb_3__1__17_chanx_right_out;
wire [0:63] sb_3__1__17_chany_bottom_out;
wire [0:63] sb_3__1__17_chany_top_out;
wire [0:63] sb_3__1__18_chanx_left_out;
wire [0:63] sb_3__1__18_chanx_right_out;
wire [0:63] sb_3__1__18_chany_bottom_out;
wire [0:63] sb_3__1__18_chany_top_out;
wire [0:0] sb_3__1__19_ccff_tail;
wire [0:63] sb_3__1__19_chanx_left_out;
wire [0:63] sb_3__1__19_chanx_right_out;
wire [0:63] sb_3__1__19_chany_bottom_out;
wire [0:63] sb_3__1__19_chany_top_out;
wire [0:0] sb_3__1__1_ccff_tail;
wire [0:63] sb_3__1__1_chanx_left_out;
wire [0:63] sb_3__1__1_chanx_right_out;
wire [0:63] sb_3__1__1_chany_bottom_out;
wire [0:63] sb_3__1__1_chany_top_out;
wire [0:0] sb_3__1__20_ccff_tail;
wire [0:63] sb_3__1__20_chanx_left_out;
wire [0:63] sb_3__1__20_chanx_right_out;
wire [0:63] sb_3__1__20_chany_bottom_out;
wire [0:63] sb_3__1__20_chany_top_out;
wire [0:0] sb_3__1__21_ccff_tail;
wire [0:63] sb_3__1__21_chanx_left_out;
wire [0:63] sb_3__1__21_chanx_right_out;
wire [0:63] sb_3__1__21_chany_bottom_out;
wire [0:63] sb_3__1__21_chany_top_out;
wire [0:0] sb_3__1__22_ccff_tail;
wire [0:63] sb_3__1__22_chanx_left_out;
wire [0:63] sb_3__1__22_chanx_right_out;
wire [0:63] sb_3__1__22_chany_bottom_out;
wire [0:63] sb_3__1__22_chany_top_out;
wire [0:0] sb_3__1__23_ccff_tail;
wire [0:63] sb_3__1__23_chanx_left_out;
wire [0:63] sb_3__1__23_chanx_right_out;
wire [0:63] sb_3__1__23_chany_bottom_out;
wire [0:63] sb_3__1__23_chany_top_out;
wire [0:0] sb_3__1__24_ccff_tail;
wire [0:63] sb_3__1__24_chanx_left_out;
wire [0:63] sb_3__1__24_chanx_right_out;
wire [0:63] sb_3__1__24_chany_bottom_out;
wire [0:63] sb_3__1__24_chany_top_out;
wire [0:0] sb_3__1__25_ccff_tail;
wire [0:63] sb_3__1__25_chanx_left_out;
wire [0:63] sb_3__1__25_chanx_right_out;
wire [0:63] sb_3__1__25_chany_bottom_out;
wire [0:63] sb_3__1__25_chany_top_out;
wire [0:0] sb_3__1__26_ccff_tail;
wire [0:63] sb_3__1__26_chanx_left_out;
wire [0:63] sb_3__1__26_chanx_right_out;
wire [0:63] sb_3__1__26_chany_bottom_out;
wire [0:63] sb_3__1__26_chany_top_out;
wire [0:0] sb_3__1__27_ccff_tail;
wire [0:63] sb_3__1__27_chanx_left_out;
wire [0:63] sb_3__1__27_chanx_right_out;
wire [0:63] sb_3__1__27_chany_bottom_out;
wire [0:63] sb_3__1__27_chany_top_out;
wire [0:0] sb_3__1__28_ccff_tail;
wire [0:63] sb_3__1__28_chanx_left_out;
wire [0:63] sb_3__1__28_chanx_right_out;
wire [0:63] sb_3__1__28_chany_bottom_out;
wire [0:63] sb_3__1__28_chany_top_out;
wire [0:0] sb_3__1__29_ccff_tail;
wire [0:63] sb_3__1__29_chanx_left_out;
wire [0:63] sb_3__1__29_chanx_right_out;
wire [0:63] sb_3__1__29_chany_bottom_out;
wire [0:63] sb_3__1__29_chany_top_out;
wire [0:0] sb_3__1__2_ccff_tail;
wire [0:63] sb_3__1__2_chanx_left_out;
wire [0:63] sb_3__1__2_chanx_right_out;
wire [0:63] sb_3__1__2_chany_bottom_out;
wire [0:63] sb_3__1__2_chany_top_out;
wire [0:0] sb_3__1__30_ccff_tail;
wire [0:63] sb_3__1__30_chanx_left_out;
wire [0:63] sb_3__1__30_chanx_right_out;
wire [0:63] sb_3__1__30_chany_bottom_out;
wire [0:63] sb_3__1__30_chany_top_out;
wire [0:0] sb_3__1__31_ccff_tail;
wire [0:63] sb_3__1__31_chanx_left_out;
wire [0:63] sb_3__1__31_chanx_right_out;
wire [0:63] sb_3__1__31_chany_bottom_out;
wire [0:63] sb_3__1__31_chany_top_out;
wire [0:0] sb_3__1__32_ccff_tail;
wire [0:63] sb_3__1__32_chanx_left_out;
wire [0:63] sb_3__1__32_chanx_right_out;
wire [0:63] sb_3__1__32_chany_bottom_out;
wire [0:63] sb_3__1__32_chany_top_out;
wire [0:0] sb_3__1__33_ccff_tail;
wire [0:63] sb_3__1__33_chanx_left_out;
wire [0:63] sb_3__1__33_chanx_right_out;
wire [0:63] sb_3__1__33_chany_bottom_out;
wire [0:63] sb_3__1__33_chany_top_out;
wire [0:0] sb_3__1__3_ccff_tail;
wire [0:63] sb_3__1__3_chanx_left_out;
wire [0:63] sb_3__1__3_chanx_right_out;
wire [0:63] sb_3__1__3_chany_bottom_out;
wire [0:63] sb_3__1__3_chany_top_out;
wire [0:0] sb_3__1__4_ccff_tail;
wire [0:63] sb_3__1__4_chanx_left_out;
wire [0:63] sb_3__1__4_chanx_right_out;
wire [0:63] sb_3__1__4_chany_bottom_out;
wire [0:63] sb_3__1__4_chany_top_out;
wire [0:0] sb_3__1__5_ccff_tail;
wire [0:63] sb_3__1__5_chanx_left_out;
wire [0:63] sb_3__1__5_chanx_right_out;
wire [0:63] sb_3__1__5_chany_bottom_out;
wire [0:63] sb_3__1__5_chany_top_out;
wire [0:0] sb_3__1__6_ccff_tail;
wire [0:63] sb_3__1__6_chanx_left_out;
wire [0:63] sb_3__1__6_chanx_right_out;
wire [0:63] sb_3__1__6_chany_bottom_out;
wire [0:63] sb_3__1__6_chany_top_out;
wire [0:0] sb_3__1__7_ccff_tail;
wire [0:63] sb_3__1__7_chanx_left_out;
wire [0:63] sb_3__1__7_chanx_right_out;
wire [0:63] sb_3__1__7_chany_bottom_out;
wire [0:63] sb_3__1__7_chany_top_out;
wire [0:0] sb_3__1__8_ccff_tail;
wire [0:63] sb_3__1__8_chanx_left_out;
wire [0:63] sb_3__1__8_chanx_right_out;
wire [0:63] sb_3__1__8_chany_bottom_out;
wire [0:63] sb_3__1__8_chany_top_out;
wire [0:0] sb_3__1__9_ccff_tail;
wire [0:63] sb_3__1__9_chanx_left_out;
wire [0:63] sb_3__1__9_chanx_right_out;
wire [0:63] sb_3__1__9_chany_bottom_out;
wire [0:63] sb_3__1__9_chany_top_out;
wire [0:0] sb_4__0__0_ccff_tail;
wire [0:63] sb_4__0__0_chanx_left_out;
wire [0:63] sb_4__0__0_chanx_right_out;
wire [0:63] sb_4__0__0_chany_top_out;
wire [0:0] sb_4__0__1_ccff_tail;
wire [0:63] sb_4__0__1_chanx_left_out;
wire [0:63] sb_4__0__1_chanx_right_out;
wire [0:63] sb_4__0__1_chany_top_out;
wire [0:0] sb_4__18__0_ccff_tail;
wire [0:63] sb_4__18__0_chanx_left_out;
wire [0:63] sb_4__18__0_chanx_right_out;
wire [0:63] sb_4__18__0_chany_bottom_out;
wire [0:0] sb_4__18__1_ccff_tail;
wire [0:63] sb_4__18__1_chanx_left_out;
wire [0:63] sb_4__18__1_chanx_right_out;
wire [0:63] sb_4__18__1_chany_bottom_out;
wire [0:0] sb_4__1__0_ccff_tail;
wire [0:63] sb_4__1__0_chanx_left_out;
wire [0:63] sb_4__1__0_chanx_right_out;
wire [0:63] sb_4__1__0_chany_bottom_out;
wire [0:63] sb_4__1__0_chany_top_out;
wire [0:0] sb_4__1__10_ccff_tail;
wire [0:63] sb_4__1__10_chanx_left_out;
wire [0:63] sb_4__1__10_chanx_right_out;
wire [0:63] sb_4__1__10_chany_bottom_out;
wire [0:63] sb_4__1__10_chany_top_out;
wire [0:0] sb_4__1__11_ccff_tail;
wire [0:63] sb_4__1__11_chanx_left_out;
wire [0:63] sb_4__1__11_chanx_right_out;
wire [0:63] sb_4__1__11_chany_bottom_out;
wire [0:63] sb_4__1__11_chany_top_out;
wire [0:0] sb_4__1__12_ccff_tail;
wire [0:63] sb_4__1__12_chanx_left_out;
wire [0:63] sb_4__1__12_chanx_right_out;
wire [0:63] sb_4__1__12_chany_bottom_out;
wire [0:63] sb_4__1__12_chany_top_out;
wire [0:0] sb_4__1__13_ccff_tail;
wire [0:63] sb_4__1__13_chanx_left_out;
wire [0:63] sb_4__1__13_chanx_right_out;
wire [0:63] sb_4__1__13_chany_bottom_out;
wire [0:63] sb_4__1__13_chany_top_out;
wire [0:0] sb_4__1__14_ccff_tail;
wire [0:63] sb_4__1__14_chanx_left_out;
wire [0:63] sb_4__1__14_chanx_right_out;
wire [0:63] sb_4__1__14_chany_bottom_out;
wire [0:63] sb_4__1__14_chany_top_out;
wire [0:0] sb_4__1__15_ccff_tail;
wire [0:63] sb_4__1__15_chanx_left_out;
wire [0:63] sb_4__1__15_chanx_right_out;
wire [0:63] sb_4__1__15_chany_bottom_out;
wire [0:63] sb_4__1__15_chany_top_out;
wire [0:0] sb_4__1__16_ccff_tail;
wire [0:63] sb_4__1__16_chanx_left_out;
wire [0:63] sb_4__1__16_chanx_right_out;
wire [0:63] sb_4__1__16_chany_bottom_out;
wire [0:63] sb_4__1__16_chany_top_out;
wire [0:0] sb_4__1__17_ccff_tail;
wire [0:63] sb_4__1__17_chanx_left_out;
wire [0:63] sb_4__1__17_chanx_right_out;
wire [0:63] sb_4__1__17_chany_bottom_out;
wire [0:63] sb_4__1__17_chany_top_out;
wire [0:0] sb_4__1__18_ccff_tail;
wire [0:63] sb_4__1__18_chanx_left_out;
wire [0:63] sb_4__1__18_chanx_right_out;
wire [0:63] sb_4__1__18_chany_bottom_out;
wire [0:63] sb_4__1__18_chany_top_out;
wire [0:0] sb_4__1__19_ccff_tail;
wire [0:63] sb_4__1__19_chanx_left_out;
wire [0:63] sb_4__1__19_chanx_right_out;
wire [0:63] sb_4__1__19_chany_bottom_out;
wire [0:63] sb_4__1__19_chany_top_out;
wire [0:0] sb_4__1__1_ccff_tail;
wire [0:63] sb_4__1__1_chanx_left_out;
wire [0:63] sb_4__1__1_chanx_right_out;
wire [0:63] sb_4__1__1_chany_bottom_out;
wire [0:63] sb_4__1__1_chany_top_out;
wire [0:0] sb_4__1__20_ccff_tail;
wire [0:63] sb_4__1__20_chanx_left_out;
wire [0:63] sb_4__1__20_chanx_right_out;
wire [0:63] sb_4__1__20_chany_bottom_out;
wire [0:63] sb_4__1__20_chany_top_out;
wire [0:0] sb_4__1__21_ccff_tail;
wire [0:63] sb_4__1__21_chanx_left_out;
wire [0:63] sb_4__1__21_chanx_right_out;
wire [0:63] sb_4__1__21_chany_bottom_out;
wire [0:63] sb_4__1__21_chany_top_out;
wire [0:0] sb_4__1__22_ccff_tail;
wire [0:63] sb_4__1__22_chanx_left_out;
wire [0:63] sb_4__1__22_chanx_right_out;
wire [0:63] sb_4__1__22_chany_bottom_out;
wire [0:63] sb_4__1__22_chany_top_out;
wire [0:0] sb_4__1__23_ccff_tail;
wire [0:63] sb_4__1__23_chanx_left_out;
wire [0:63] sb_4__1__23_chanx_right_out;
wire [0:63] sb_4__1__23_chany_bottom_out;
wire [0:63] sb_4__1__23_chany_top_out;
wire [0:0] sb_4__1__24_ccff_tail;
wire [0:63] sb_4__1__24_chanx_left_out;
wire [0:63] sb_4__1__24_chanx_right_out;
wire [0:63] sb_4__1__24_chany_bottom_out;
wire [0:63] sb_4__1__24_chany_top_out;
wire [0:0] sb_4__1__25_ccff_tail;
wire [0:63] sb_4__1__25_chanx_left_out;
wire [0:63] sb_4__1__25_chanx_right_out;
wire [0:63] sb_4__1__25_chany_bottom_out;
wire [0:63] sb_4__1__25_chany_top_out;
wire [0:0] sb_4__1__26_ccff_tail;
wire [0:63] sb_4__1__26_chanx_left_out;
wire [0:63] sb_4__1__26_chanx_right_out;
wire [0:63] sb_4__1__26_chany_bottom_out;
wire [0:63] sb_4__1__26_chany_top_out;
wire [0:0] sb_4__1__27_ccff_tail;
wire [0:63] sb_4__1__27_chanx_left_out;
wire [0:63] sb_4__1__27_chanx_right_out;
wire [0:63] sb_4__1__27_chany_bottom_out;
wire [0:63] sb_4__1__27_chany_top_out;
wire [0:0] sb_4__1__28_ccff_tail;
wire [0:63] sb_4__1__28_chanx_left_out;
wire [0:63] sb_4__1__28_chanx_right_out;
wire [0:63] sb_4__1__28_chany_bottom_out;
wire [0:63] sb_4__1__28_chany_top_out;
wire [0:0] sb_4__1__29_ccff_tail;
wire [0:63] sb_4__1__29_chanx_left_out;
wire [0:63] sb_4__1__29_chanx_right_out;
wire [0:63] sb_4__1__29_chany_bottom_out;
wire [0:63] sb_4__1__29_chany_top_out;
wire [0:0] sb_4__1__2_ccff_tail;
wire [0:63] sb_4__1__2_chanx_left_out;
wire [0:63] sb_4__1__2_chanx_right_out;
wire [0:63] sb_4__1__2_chany_bottom_out;
wire [0:63] sb_4__1__2_chany_top_out;
wire [0:0] sb_4__1__30_ccff_tail;
wire [0:63] sb_4__1__30_chanx_left_out;
wire [0:63] sb_4__1__30_chanx_right_out;
wire [0:63] sb_4__1__30_chany_bottom_out;
wire [0:63] sb_4__1__30_chany_top_out;
wire [0:0] sb_4__1__31_ccff_tail;
wire [0:63] sb_4__1__31_chanx_left_out;
wire [0:63] sb_4__1__31_chanx_right_out;
wire [0:63] sb_4__1__31_chany_bottom_out;
wire [0:63] sb_4__1__31_chany_top_out;
wire [0:0] sb_4__1__32_ccff_tail;
wire [0:63] sb_4__1__32_chanx_left_out;
wire [0:63] sb_4__1__32_chanx_right_out;
wire [0:63] sb_4__1__32_chany_bottom_out;
wire [0:63] sb_4__1__32_chany_top_out;
wire [0:0] sb_4__1__33_ccff_tail;
wire [0:63] sb_4__1__33_chanx_left_out;
wire [0:63] sb_4__1__33_chanx_right_out;
wire [0:63] sb_4__1__33_chany_bottom_out;
wire [0:63] sb_4__1__33_chany_top_out;
wire [0:0] sb_4__1__3_ccff_tail;
wire [0:63] sb_4__1__3_chanx_left_out;
wire [0:63] sb_4__1__3_chanx_right_out;
wire [0:63] sb_4__1__3_chany_bottom_out;
wire [0:63] sb_4__1__3_chany_top_out;
wire [0:0] sb_4__1__4_ccff_tail;
wire [0:63] sb_4__1__4_chanx_left_out;
wire [0:63] sb_4__1__4_chanx_right_out;
wire [0:63] sb_4__1__4_chany_bottom_out;
wire [0:63] sb_4__1__4_chany_top_out;
wire [0:0] sb_4__1__5_ccff_tail;
wire [0:63] sb_4__1__5_chanx_left_out;
wire [0:63] sb_4__1__5_chanx_right_out;
wire [0:63] sb_4__1__5_chany_bottom_out;
wire [0:63] sb_4__1__5_chany_top_out;
wire [0:0] sb_4__1__6_ccff_tail;
wire [0:63] sb_4__1__6_chanx_left_out;
wire [0:63] sb_4__1__6_chanx_right_out;
wire [0:63] sb_4__1__6_chany_bottom_out;
wire [0:63] sb_4__1__6_chany_top_out;
wire [0:0] sb_4__1__7_ccff_tail;
wire [0:63] sb_4__1__7_chanx_left_out;
wire [0:63] sb_4__1__7_chanx_right_out;
wire [0:63] sb_4__1__7_chany_bottom_out;
wire [0:63] sb_4__1__7_chany_top_out;
wire [0:0] sb_4__1__8_ccff_tail;
wire [0:63] sb_4__1__8_chanx_left_out;
wire [0:63] sb_4__1__8_chanx_right_out;
wire [0:63] sb_4__1__8_chany_bottom_out;
wire [0:63] sb_4__1__8_chany_top_out;
wire [0:0] sb_4__1__9_ccff_tail;
wire [0:63] sb_4__1__9_chanx_left_out;
wire [0:63] sb_4__1__9_chanx_right_out;
wire [0:63] sb_4__1__9_chany_bottom_out;
wire [0:63] sb_4__1__9_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_clb grid_clb_1__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_204_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_205_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_206_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_207_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_208_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_1__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_209_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_1__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_210_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_1__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_211_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_1__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_212_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_1__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_213_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_1__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_214_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_1__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_215_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_1__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_216_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_1__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_217_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_1__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_218_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_1__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_219_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_1__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_220_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_1__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__18__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail[11]));

	grid_clb grid_clb_2__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_221_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_222_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_223_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_224_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_225_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__22_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_2__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_226_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__23_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_2__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_227_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__24_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_24_ccff_tail));

	grid_clb grid_clb_2__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_228_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__25_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_25_ccff_tail));

	grid_clb grid_clb_2__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_229_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__26_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_26_ccff_tail));

	grid_clb grid_clb_2__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_230_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__27_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_27_ccff_tail));

	grid_clb grid_clb_2__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_231_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__28_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_28_ccff_tail));

	grid_clb grid_clb_2__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_232_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_28_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__29_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_29_ccff_tail));

	grid_clb grid_clb_2__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_233_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_29_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__30_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_30_ccff_tail));

	grid_clb grid_clb_2__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_234_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_30_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__31_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_31_ccff_tail));

	grid_clb grid_clb_2__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_235_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_31_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__32_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_32_ccff_tail));

	grid_clb grid_clb_2__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_236_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_32_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__33_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_33_ccff_tail));

	grid_clb grid_clb_2__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_237_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_33_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__34_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail[10]));

	grid_clb grid_clb_2__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_408_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__35_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_35_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_238_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_34_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_36_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_239_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_35_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_37_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_240_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_36_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_38_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_241_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_37_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_39_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_242_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_38_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_40_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_243_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_39_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_41_ccff_tail));

	grid_clb grid_clb_3__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_244_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_40_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_42_ccff_tail));

	grid_clb grid_clb_3__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_245_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_41_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_43_ccff_tail));

	grid_clb grid_clb_3__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_246_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_42_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_44_ccff_tail));

	grid_clb grid_clb_3__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_247_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_43_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_45_ccff_tail));

	grid_clb grid_clb_3__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_248_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_44_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_46_ccff_tail));

	grid_clb grid_clb_3__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_249_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_45_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_47_ccff_tail));

	grid_clb grid_clb_3__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_250_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_46_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_48_ccff_tail));

	grid_clb grid_clb_3__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_251_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_47_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_49_ccff_tail));

	grid_clb grid_clb_3__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_252_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_48_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_50_ccff_tail));

	grid_clb grid_clb_3__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_253_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_49_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_51_ccff_tail));

	grid_clb grid_clb_3__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_254_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_50_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_52_ccff_tail));

	grid_clb grid_clb_3__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_409_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_53_ccff_tail));

	grid_clb grid_clb_5__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_255_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_51_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__36_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_54_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_256_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_52_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__37_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_55_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_257_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_53_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__38_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_56_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_258_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_54_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__39_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_57_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_259_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_55_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__40_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail[3]));

	grid_clb grid_clb_5__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_260_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_56_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__41_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_59_ccff_tail));

	grid_clb grid_clb_5__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_261_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_57_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__42_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_60_ccff_tail));

	grid_clb grid_clb_5__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_262_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_58_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__43_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail[5]));

	grid_clb grid_clb_5__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_263_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_59_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__44_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_62_ccff_tail));

	grid_clb grid_clb_5__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_264_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_60_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__45_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_63_ccff_tail));

	grid_clb grid_clb_5__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_265_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_61_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__46_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_64_ccff_tail));

	grid_clb grid_clb_5__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_266_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_62_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__47_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_65_ccff_tail));

	grid_clb grid_clb_5__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_267_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_63_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__48_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_66_ccff_tail));

	grid_clb grid_clb_5__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_268_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_64_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__49_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_67_ccff_tail));

	grid_clb grid_clb_5__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_269_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_65_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__50_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_68_ccff_tail));

	grid_clb grid_clb_5__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_270_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_66_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__51_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_69_ccff_tail));

	grid_clb grid_clb_5__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_271_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_67_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__52_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_70_ccff_tail));

	grid_clb grid_clb_5__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_410_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__53_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_71_ccff_tail));

	grid_clb grid_clb_6__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_272_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_68_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__54_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_72_ccff_tail));

	grid_clb grid_clb_6__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_273_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_69_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__55_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_73_ccff_tail));

	grid_clb grid_clb_6__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_274_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_70_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__56_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_74_ccff_tail));

	grid_clb grid_clb_6__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_275_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_71_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__57_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_75_ccff_tail));

	grid_clb grid_clb_6__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_276_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_72_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__58_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_76_ccff_tail));

	grid_clb grid_clb_6__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_277_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_73_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__59_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_77_ccff_tail));

	grid_clb grid_clb_6__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_278_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_74_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__60_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_78_ccff_tail));

	grid_clb grid_clb_6__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_279_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_75_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__61_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_79_ccff_tail));

	grid_clb grid_clb_6__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_280_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_76_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__62_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_80_ccff_tail));

	grid_clb grid_clb_6__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_281_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_77_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__63_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_81_ccff_tail));

	grid_clb grid_clb_6__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_282_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_78_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__64_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_82_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_82_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_82_ccff_tail));

	grid_clb grid_clb_6__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_283_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_79_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__65_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_83_ccff_tail));

	grid_clb grid_clb_6__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_284_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_80_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__66_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_84_ccff_tail));

	grid_clb grid_clb_6__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_285_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_81_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__67_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_85_ccff_tail));

	grid_clb grid_clb_6__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_286_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_82_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__68_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_86_ccff_tail));

	grid_clb grid_clb_6__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_287_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_83_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__69_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_87_ccff_tail));

	grid_clb grid_clb_6__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_288_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_84_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__70_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_88_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_88_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_88_ccff_tail));

	grid_clb grid_clb_6__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_411_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__71_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_89_ccff_tail));

	grid_clb grid_clb_7__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_289_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_85_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__72_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_90_ccff_tail));

	grid_clb grid_clb_7__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_290_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_86_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__73_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_91_ccff_tail));

	grid_clb grid_clb_7__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_291_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_87_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__74_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_92_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_92_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_92_ccff_tail));

	grid_clb grid_clb_7__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_292_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_88_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__75_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_93_ccff_tail));

	grid_clb grid_clb_7__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_293_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_89_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__76_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_94_ccff_tail));

	grid_clb grid_clb_7__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_294_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_90_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__77_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_95_ccff_tail));

	grid_clb grid_clb_7__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_295_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_91_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__78_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_96_ccff_tail));

	grid_clb grid_clb_7__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_296_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_92_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__79_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_97_ccff_tail));

	grid_clb grid_clb_7__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_297_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_93_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__80_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_98_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_98_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_98_ccff_tail));

	grid_clb grid_clb_7__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_298_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_94_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__81_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_99_ccff_tail));

	grid_clb grid_clb_7__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_299_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_95_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__82_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_100_ccff_tail));

	grid_clb grid_clb_7__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_300_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_96_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__83_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_101_ccff_tail));

	grid_clb grid_clb_7__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_301_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_97_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__84_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_102_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_102_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_102_ccff_tail));

	grid_clb grid_clb_7__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_302_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_98_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__85_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_103_ccff_tail));

	grid_clb grid_clb_7__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_303_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_99_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__86_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_104_ccff_tail));

	grid_clb grid_clb_7__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_304_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_100_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__87_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_105_ccff_tail));

	grid_clb grid_clb_7__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_305_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_101_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__88_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_106_ccff_tail));

	grid_clb grid_clb_7__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_412_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__89_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_107_ccff_tail));

	grid_clb grid_clb_8__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_306_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_102_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__90_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_108_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_108_ccff_tail));

	grid_clb grid_clb_8__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_307_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_103_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__91_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_109_ccff_tail));

	grid_clb grid_clb_8__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_308_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_104_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__92_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_110_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_110_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_110_ccff_tail));

	grid_clb grid_clb_8__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_309_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_105_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__93_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_111_ccff_tail));

	grid_clb grid_clb_8__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_310_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_106_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__94_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_112_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_112_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_112_ccff_tail));

	grid_clb grid_clb_8__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_311_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_107_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__95_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_113_ccff_tail));

	grid_clb grid_clb_8__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_312_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_108_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__96_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_114_ccff_tail));

	grid_clb grid_clb_8__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_313_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_109_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__97_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_115_ccff_tail));

	grid_clb grid_clb_8__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_314_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_110_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__98_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_116_ccff_tail));

	grid_clb grid_clb_8__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_315_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_111_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__99_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_117_ccff_tail));

	grid_clb grid_clb_8__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_316_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_112_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__100_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_118_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_118_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_118_ccff_tail));

	grid_clb grid_clb_8__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_317_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_113_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__101_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_119_ccff_tail));

	grid_clb grid_clb_8__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_318_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_114_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__102_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_120_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_120_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_120_ccff_tail));

	grid_clb grid_clb_8__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_319_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_115_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__103_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_121_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_121_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_121_ccff_tail));

	grid_clb grid_clb_8__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_320_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_116_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__104_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_122_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_122_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_122_ccff_tail));

	grid_clb grid_clb_8__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_321_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_117_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__105_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_123_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_123_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_123_ccff_tail));

	grid_clb grid_clb_8__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_322_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_118_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__106_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_124_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_124_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_124_ccff_tail));

	grid_clb grid_clb_8__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_413_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__107_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_125_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_125_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_125_ccff_tail));

	grid_clb grid_clb_9__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_323_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_119_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__108_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_126_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_126_ccff_tail));

	grid_clb grid_clb_9__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_324_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_120_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__109_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_127_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_127_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_127_ccff_tail));

	grid_clb grid_clb_9__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_325_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_121_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__110_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_128_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_128_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_128_ccff_tail));

	grid_clb grid_clb_9__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_326_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_122_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__111_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_129_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_129_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_129_ccff_tail));

	grid_clb grid_clb_9__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_327_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_123_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__112_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_130_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_130_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_130_ccff_tail));

	grid_clb grid_clb_9__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_328_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_124_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__113_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_131_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_131_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_131_ccff_tail));

	grid_clb grid_clb_9__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_329_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_125_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__114_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_132_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_132_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_132_ccff_tail));

	grid_clb grid_clb_9__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_330_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_126_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__115_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_133_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_133_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_133_ccff_tail));

	grid_clb grid_clb_9__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_331_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_127_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__116_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_134_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_134_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_134_ccff_tail));

	grid_clb grid_clb_9__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_332_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_128_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(ccff_head[7]),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_135_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_135_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_135_ccff_tail));

	grid_clb grid_clb_9__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_333_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_129_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__118_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_136_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_136_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_136_ccff_tail));

	grid_clb grid_clb_9__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_334_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_130_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__119_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_137_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_137_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_137_ccff_tail));

	grid_clb grid_clb_9__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_335_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_131_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__120_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_138_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_138_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_138_ccff_tail));

	grid_clb grid_clb_9__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_336_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_132_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__121_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_139_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_139_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_139_ccff_tail));

	grid_clb grid_clb_9__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_337_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_133_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__122_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_140_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_140_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_140_ccff_tail));

	grid_clb grid_clb_9__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_338_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_134_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__123_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_141_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_141_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_141_ccff_tail));

	grid_clb grid_clb_9__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_339_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_135_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__124_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_142_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_142_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_142_ccff_tail));

	grid_clb grid_clb_9__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_414_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__125_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_143_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_143_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_143_ccff_tail));

	grid_clb grid_clb_10__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_340_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_136_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_144_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_144_ccff_tail));

	grid_clb grid_clb_10__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_341_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_137_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_145_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_145_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_145_ccff_tail));

	grid_clb grid_clb_10__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_342_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_138_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_146_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_146_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_146_ccff_tail));

	grid_clb grid_clb_10__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_343_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_139_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_147_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_147_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_147_ccff_tail));

	grid_clb grid_clb_10__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_344_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_140_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_148_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_148_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_148_ccff_tail));

	grid_clb grid_clb_10__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_345_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_141_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_149_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_149_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_149_ccff_tail));

	grid_clb grid_clb_10__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_346_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_142_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_150_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_150_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_150_ccff_tail));

	grid_clb grid_clb_10__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_347_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_143_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_151_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_151_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_151_ccff_tail));

	grid_clb grid_clb_10__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_348_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_144_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_152_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_152_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_152_ccff_tail));

	grid_clb grid_clb_10__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_349_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_145_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_153_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_153_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_153_ccff_tail));

	grid_clb grid_clb_10__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_350_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_146_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_154_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_154_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_154_ccff_tail));

	grid_clb grid_clb_10__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_351_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_147_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_155_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_155_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_155_ccff_tail));

	grid_clb grid_clb_10__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_352_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_148_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_156_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_156_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_156_ccff_tail));

	grid_clb grid_clb_10__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_353_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_149_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_157_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_157_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_157_ccff_tail));

	grid_clb grid_clb_10__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_354_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_150_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_158_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_158_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_158_ccff_tail));

	grid_clb grid_clb_10__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_355_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_151_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_159_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_159_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_159_ccff_tail));

	grid_clb grid_clb_10__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_356_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_152_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_160_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_160_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_160_ccff_tail));

	grid_clb grid_clb_10__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_415_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_10__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_3__2__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_161_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_161_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_161_ccff_tail));

	grid_clb grid_clb_12__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_357_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_153_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__126_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_162_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_162_ccff_tail));

	grid_clb grid_clb_12__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_358_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_154_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__127_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_163_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_163_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_163_ccff_tail));

	grid_clb grid_clb_12__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_359_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_155_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__128_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_164_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_164_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_164_ccff_tail));

	grid_clb grid_clb_12__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_360_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_156_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__129_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_165_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_165_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_165_ccff_tail));

	grid_clb grid_clb_12__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_361_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_157_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__130_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_166_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_166_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_166_ccff_tail));

	grid_clb grid_clb_12__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_362_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_158_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__131_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_167_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_167_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_167_ccff_tail));

	grid_clb grid_clb_12__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_363_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_159_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__132_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_168_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_168_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_168_ccff_tail));

	grid_clb grid_clb_12__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_364_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_160_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__133_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_169_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_169_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_169_ccff_tail));

	grid_clb grid_clb_12__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_365_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_161_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__134_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_170_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_170_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_170_ccff_tail));

	grid_clb grid_clb_12__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_366_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_162_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__135_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_171_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_171_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_171_ccff_tail));

	grid_clb grid_clb_12__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_367_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_163_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__136_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_172_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_172_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_172_ccff_tail));

	grid_clb grid_clb_12__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_368_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_164_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__137_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_173_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_173_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_173_ccff_tail));

	grid_clb grid_clb_12__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_369_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_165_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__138_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_174_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_174_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_174_ccff_tail));

	grid_clb grid_clb_12__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_370_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_166_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__139_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_175_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_175_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_175_ccff_tail));

	grid_clb grid_clb_12__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_371_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_167_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__140_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_176_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_176_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_176_ccff_tail));

	grid_clb grid_clb_12__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_372_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_168_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__141_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_177_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_177_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_177_ccff_tail));

	grid_clb grid_clb_12__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_373_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_169_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__142_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_178_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_178_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_178_ccff_tail));

	grid_clb grid_clb_12__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_416_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_12__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__143_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_179_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_179_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_179_ccff_tail));

	grid_clb grid_clb_13__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_374_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_170_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__144_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_180_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_180_ccff_tail));

	grid_clb grid_clb_13__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_375_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_171_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__145_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_181_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_181_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_181_ccff_tail));

	grid_clb grid_clb_13__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_376_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_172_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__146_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_182_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_182_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_182_ccff_tail));

	grid_clb grid_clb_13__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_377_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_173_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__147_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_183_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_183_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_183_ccff_tail));

	grid_clb grid_clb_13__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_378_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_174_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__148_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_184_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_184_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_184_ccff_tail));

	grid_clb grid_clb_13__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_379_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_175_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__149_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_185_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_185_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_185_ccff_tail));

	grid_clb grid_clb_13__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_380_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_176_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__150_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_186_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_186_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_186_ccff_tail));

	grid_clb grid_clb_13__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_381_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_177_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__151_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_187_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_187_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_187_ccff_tail));

	grid_clb grid_clb_13__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_382_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_178_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__152_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_188_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_188_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_188_ccff_tail));

	grid_clb grid_clb_13__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_383_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_179_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__153_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_189_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_189_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_189_ccff_tail));

	grid_clb grid_clb_13__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_384_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_180_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__154_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_190_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_190_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_190_ccff_tail));

	grid_clb grid_clb_13__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_385_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_181_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__155_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_191_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_191_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_191_ccff_tail));

	grid_clb grid_clb_13__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_386_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_182_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__156_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_192_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_192_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_192_ccff_tail));

	grid_clb grid_clb_13__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_387_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_183_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__157_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_193_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_193_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_193_ccff_tail));

	grid_clb grid_clb_13__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_388_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_184_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__158_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_194_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_194_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_194_ccff_tail));

	grid_clb grid_clb_13__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_389_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_185_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__159_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_195_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_195_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_195_ccff_tail));

	grid_clb grid_clb_13__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_390_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_186_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__160_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_196_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_196_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_196_ccff_tail));

	grid_clb grid_clb_13__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_417_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_13__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__161_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_197_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_197_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_197_ccff_tail));

	grid_clb grid_clb_14__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_391_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_187_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(ccff_head[2]),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_198_ccff_tail));

	grid_clb grid_clb_14__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_392_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_188_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_199_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_199_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_199_ccff_tail));

	grid_clb grid_clb_14__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_393_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_189_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_200_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_200_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_200_ccff_tail));

	grid_clb grid_clb_14__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_394_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_190_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_201_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_201_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_201_ccff_tail));

	grid_clb grid_clb_14__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_395_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_191_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_202_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_202_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_202_ccff_tail));

	grid_clb grid_clb_14__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_396_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_192_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_203_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_203_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_203_ccff_tail));

	grid_clb grid_clb_14__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_397_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_193_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_204_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_204_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_204_ccff_tail));

	grid_clb grid_clb_14__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_398_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_194_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_205_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_205_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_205_ccff_tail));

	grid_clb grid_clb_14__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_399_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_195_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_206_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_206_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_206_ccff_tail));

	grid_clb grid_clb_14__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_400_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_196_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_207_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_207_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_207_ccff_tail));

	grid_clb grid_clb_14__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_401_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_197_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_208_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_208_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_208_ccff_tail));

	grid_clb grid_clb_14__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_402_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_198_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_209_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_209_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_209_ccff_tail));

	grid_clb grid_clb_14__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_403_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_199_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_210_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_210_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_210_ccff_tail));

	grid_clb grid_clb_14__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_404_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_200_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_211_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_211_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_211_ccff_tail));

	grid_clb grid_clb_14__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_405_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_201_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_212_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_212_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_212_ccff_tail));

	grid_clb grid_clb_14__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_406_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_202_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_213_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_213_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_213_ccff_tail));

	grid_clb grid_clb_14__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_407_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_203_out),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_214_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_214_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_214_ccff_tail));

	grid_clb grid_clb_14__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_418_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_14__18__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_14__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.right_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.right_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_215_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_215_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_215_ccff_tail));

	grid_memory grid_memory_4__1_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__3_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__5_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__7_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__9_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__11_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__13_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__13__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__15_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__15__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_4__17_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_4__17__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__1_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__3_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__5_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__7_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__9_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__11_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__13_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__13__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__15_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__15__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_memory grid_memory_11__17_ (
		.top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.right_width_0_height_1_subtile_0__pin_waddr_3_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_1_subtile_0__pin_raddr_2_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_1_subtile_0__pin_data_in_1_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_1_subtile_0__pin_ren_0_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_11__17__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.top_width_0_height_0_subtile_0__pin_data_out_4_upper(grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.top_width_0_height_0_subtile_0__pin_data_out_4_lower(grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.top_width_0_height_1_subtile_0__pin_data_out_5_upper(grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.top_width_0_height_1_subtile_0__pin_data_out_5_lower(grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.right_width_0_height_0_subtile_0__pin_data_out_6_upper(grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.right_width_0_height_0_subtile_0__pin_data_out_6_lower(grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.right_width_0_height_1_subtile_0__pin_data_out_7_upper(grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.right_width_0_height_1_subtile_0__pin_data_out_7_lower(grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_upper(grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_data_out_0_lower(grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_upper(grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.bottom_width_0_height_1_subtile_0__pin_data_out_1_lower(grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_width_0_height_0_subtile_0__pin_data_out_2_upper(grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.left_width_0_height_0_subtile_0__pin_data_out_2_lower(grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.left_width_0_height_1_subtile_0__pin_data_out_3_upper(grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.left_width_0_height_1_subtile_0__pin_data_out_3_lower(grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_lower));

	grid_io_top_top grid_io_top_top_1__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[0]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[0]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[0]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_0_ccff_tail));

	grid_io_top_top grid_io_top_top_2__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[1]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[1]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[1]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_1_ccff_tail));

	grid_io_top_top grid_io_top_top_3__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[2]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[2]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[2]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_2_ccff_tail));

	grid_io_top_top grid_io_top_top_4__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[3]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[3]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[3]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_4__18__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_3_ccff_tail));

	grid_io_top_top grid_io_top_top_5__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[4]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[4]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[4]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_4_ccff_tail));

	grid_io_top_top grid_io_top_top_6__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[5]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[5]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[5]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_5_ccff_tail));

	grid_io_top_top grid_io_top_top_7__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[6]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[6]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[6]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_6_ccff_tail));

	grid_io_top_top grid_io_top_top_8__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[7]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[7]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__6_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_7_ccff_tail));

	grid_io_top_top grid_io_top_top_9__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[8]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[8]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[8]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__7_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_8_ccff_tail));

	grid_io_top_top grid_io_top_top_10__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[9]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[9]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[9]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__8_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_9_ccff_tail));

	grid_io_top_top grid_io_top_top_11__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[10]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[10]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[10]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_4__18__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_10_ccff_tail));

	grid_io_top_top grid_io_top_top_12__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[11]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[11]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[11]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__9_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_11_ccff_tail));

	grid_io_top_top grid_io_top_top_13__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[12]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[12]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[12]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__10_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_12_ccff_tail));

	grid_io_top_top grid_io_top_top_14__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[13]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[13]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[13]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__18__11_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_13_ccff_tail));

	grid_io_right_right grid_io_right_right_15__18_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[14]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[14]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[14]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_0_ccff_tail));

	grid_io_right_right grid_io_right_right_15__17_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[15]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[15]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[15]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_1_ccff_tail));

	grid_io_right_right grid_io_right_right_15__16_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[16]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[16]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[16]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_2_ccff_tail));

	grid_io_right_right grid_io_right_right_15__15_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[17]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[17]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[17]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_3_ccff_tail));

	grid_io_right_right grid_io_right_right_15__14_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[18]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[18]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[18]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_4_ccff_tail));

	grid_io_right_right grid_io_right_right_15__13_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[19]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[19]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[19]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_5_ccff_tail));

	grid_io_right_right grid_io_right_right_15__12_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[20]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[20]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[20]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_6_ccff_tail));

	grid_io_right_right grid_io_right_right_15__11_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[21]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[21]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[21]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_8_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_7_ccff_tail));

	grid_io_right_right grid_io_right_right_15__10_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[22]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[22]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[22]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_9_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_8_ccff_tail));

	grid_io_right_right grid_io_right_right_15__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[23]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[23]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[23]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_10_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_9_ccff_tail));

	grid_io_right_right grid_io_right_right_15__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[24]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[24]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[24]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_11_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_10_ccff_tail));

	grid_io_right_right grid_io_right_right_15__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[25]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[25]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[25]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_12_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_11_ccff_tail));

	grid_io_right_right grid_io_right_right_15__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[26]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[26]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[26]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_13_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_12_ccff_tail));

	grid_io_right_right grid_io_right_right_15__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[27]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[27]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[27]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_14_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_13_ccff_tail));

	grid_io_right_right grid_io_right_right_15__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[28]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[28]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[28]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_15_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_14_ccff_tail));

	grid_io_right_right grid_io_right_right_15__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[29]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[29]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[29]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_16_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_15_ccff_tail));

	grid_io_right_right grid_io_right_right_15__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[30]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[30]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[30]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_17_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_16_ccff_tail));

	grid_io_right_right grid_io_right_right_15__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[31]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[31]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[31]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_17_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_14__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[32:40]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[32:40]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[32:40]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_0_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_13__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[41:49]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[41:49]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[41:49]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_1_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_12__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[50:58]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[50:58]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[50:58]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_2_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_11__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[59:67]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[59:67]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[59:67]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_3_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_10__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[68:76]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[68:76]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[68:76]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_4_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_9__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[77:85]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[77:85]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[77:85]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_5_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_8__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[86:94]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[86:94]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[86:94]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_6_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_7__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[95:103]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[95:103]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[95:103]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_7_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_6__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[104:112]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[104:112]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[104:112]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_8_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_5__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[113:121]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[113:121]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[113:121]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_9_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_4__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[122:130]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[122:130]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[122:130]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_10_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_3__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[131:139]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[131:139]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[131:139]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_11_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_2__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[140:148]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[140:148]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[140:148]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_12_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_1__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[149:157]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[149:157]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[149:157]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(ccff_head[0]),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_13_ccff_tail));

	grid_io_left_left grid_io_left_left_0__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[158]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[158]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[158]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_0_ccff_tail));

	grid_io_left_left grid_io_left_left_0__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[159]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[159]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[159]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_1_ccff_tail));

	grid_io_left_left grid_io_left_left_0__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[160]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[160]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[160]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_2_ccff_tail));

	grid_io_left_left grid_io_left_left_0__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[161]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[161]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[161]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_3_ccff_tail));

	grid_io_left_left grid_io_left_left_0__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[162]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[162]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[162]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_4_ccff_tail));

	grid_io_left_left grid_io_left_left_0__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[163]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[163]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[163]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_5_ccff_tail));

	grid_io_left_left grid_io_left_left_0__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[164]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[164]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[164]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_6_ccff_tail));

	grid_io_left_left grid_io_left_left_0__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[165]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[165]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[165]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_7_ccff_tail));

	grid_io_left_left grid_io_left_left_0__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[166]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[166]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[166]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__8_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_8_ccff_tail));

	grid_io_left_left grid_io_left_left_0__10_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[167]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[167]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[167]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__9_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_9_ccff_tail));

	grid_io_left_left grid_io_left_left_0__11_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[168]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[168]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[168]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__10_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_10_ccff_tail));

	grid_io_left_left grid_io_left_left_0__12_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[169]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[169]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[169]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__11_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_11_ccff_tail));

	grid_io_left_left grid_io_left_left_0__13_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[170]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[170]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[170]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__12_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_12_ccff_tail));

	grid_io_left_left grid_io_left_left_0__14_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[171]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[171]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[171]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__13_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_13_ccff_tail));

	grid_io_left_left grid_io_left_left_0__15_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[172]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[172]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[172]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__14_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_14_ccff_tail));

	grid_io_left_left grid_io_left_left_0__16_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[173]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[173]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[173]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__15_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_15_ccff_tail));

	grid_io_left_left grid_io_left_left_0__17_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[174]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[174]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[174]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__16_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_16_ccff_tail));

	grid_io_left_left grid_io_left_left_0__18_ (
		.IO_ISOL_N(IO_ISOL_N),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[175]),
		.gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[175]),
		.gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[175]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__17_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_17_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:63]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:63]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_4_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_5_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__1_ sb_0__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_6_ccff_tail),
		.chany_top_out(sb_0__1__4_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__4_ccff_tail));

	sb_0__1_ sb_0__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_7_ccff_tail),
		.chany_top_out(sb_0__1__5_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__5_ccff_tail));

	sb_0__1_ sb_0__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_8_ccff_tail),
		.chany_top_out(sb_0__1__6_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__6_ccff_tail));

	sb_0__1_ sb_0__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__8_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_9_ccff_tail),
		.chany_top_out(sb_0__1__7_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__7_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__7_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__7_ccff_tail));

	sb_0__1_ sb_0__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__9_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_10_ccff_tail),
		.chany_top_out(sb_0__1__8_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__8_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__8_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__8_ccff_tail));

	sb_0__1_ sb_0__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__10_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_11_ccff_tail),
		.chany_top_out(sb_0__1__9_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__9_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__9_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__9_ccff_tail));

	sb_0__1_ sb_0__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__11_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__10_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_12_ccff_tail),
		.chany_top_out(sb_0__1__10_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__10_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__10_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__10_ccff_tail));

	sb_0__1_ sb_0__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__12_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__11_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_13_ccff_tail),
		.chany_top_out(sb_0__1__11_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__11_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__11_chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[0]));

	sb_0__1_ sb_0__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__13_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__12_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_14_ccff_tail),
		.chany_top_out(sb_0__1__12_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__12_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__12_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__12_ccff_tail));

	sb_0__1_ sb_0__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__14_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__13_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_15_ccff_tail),
		.chany_top_out(sb_0__1__13_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__13_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__13_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__13_ccff_tail));

	sb_0__1_ sb_0__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__15_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__14_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_16_ccff_tail),
		.chany_top_out(sb_0__1__14_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__14_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__14_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__14_ccff_tail));

	sb_0__1_ sb_0__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__16_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__15_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_17_ccff_tail),
		.chany_top_out(sb_0__1__15_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__15_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__15_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__15_ccff_tail));

	sb_0__1_ sb_0__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__17_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__16_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(sb_0__18__0_ccff_tail),
		.chany_top_out(sb_0__1__16_chany_top_out[0:63]),
		.chanx_right_out(sb_0__1__16_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__1__16_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__1__16_ccff_tail));

	sb_0__18_ sb_0__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__0_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_0__1__17_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_top_top_0_ccff_tail),
		.chanx_right_out(sb_0__18__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_0__18__0_chany_bottom_out[0:63]),
		.ccff_tail(sb_0__18__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__18_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_13_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_io_left_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__36_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__18_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_12_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_5__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__36_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__72_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__54_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(cby_4__1__0_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_6__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__54_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__90_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__72_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_54_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_7__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__72_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__108_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__90_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_72_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__0_ sb_8__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__90_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__126_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__108_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_90_ccff_tail),
		.chany_top_out(sb_1__0__5_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__5_ccff_tail));

	sb_1__0_ sb_9__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__108_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__144_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__126_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_108_ccff_tail),
		.chany_top_out(sb_1__0__6_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__6_ccff_tail));

	sb_1__0_ sb_12__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__126_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__180_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__162_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(cby_4__1__18_ccff_tail),
		.chany_top_out(sb_1__0__7_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__7_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__7_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__7_ccff_tail));

	sb_1__0_ sb_13__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__144_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__198_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__180_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_162_ccff_tail),
		.chany_top_out(sb_1__0__8_chany_top_out[0:63]),
		.chanx_right_out(sb_1__0__8_chanx_right_out[0:63]),
		.chanx_left_out(sb_1__0__8_chanx_left_out[0:63]),
		.ccff_tail(sb_1__0__8_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__19_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__20_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__21_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_1__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__22_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_1__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__23_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_1__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__24_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_1__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__25_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_25_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_1__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__26_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__8_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_1__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__27_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__9_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_27_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__1_ sb_1__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__28_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__10_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__1__9_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__9_ccff_tail));

	sb_1__1_ sb_1__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__29_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__11_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_29_ccff_tail),
		.chany_top_out(sb_1__1__10_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__10_ccff_tail));

	sb_1__1_ sb_1__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__30_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__12_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__1__11_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__11_ccff_tail));

	sb_1__1_ sb_1__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__31_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__13_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_31_ccff_tail),
		.chany_top_out(sb_1__1__12_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__12_ccff_tail));

	sb_1__1_ sb_1__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__32_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__14_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__1__13_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__13_ccff_tail));

	sb_1__1_ sb_1__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__33_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__15_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_33_ccff_tail),
		.chany_top_out(sb_1__1__14_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__14_ccff_tail));

	sb_1__1_ sb_1__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__34_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__16_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__1__15_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__15_ccff_tail));

	sb_1__1_ sb_1__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__35_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__17_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_35_ccff_tail),
		.chany_top_out(sb_1__1__16_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__16_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__37_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__19_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_37_ccff_tail),
		.chany_top_out(sb_1__1__17_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__17_ccff_tail));

	sb_1__1_ sb_2__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__20_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__38_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__20_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__18_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__18_ccff_tail));

	sb_1__1_ sb_2__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__21_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__39_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__21_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_39_ccff_tail),
		.chany_top_out(sb_1__1__19_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__19_ccff_tail));

	sb_1__1_ sb_2__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__22_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__40_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__22_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__1__20_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__20_ccff_tail));

	sb_1__1_ sb_2__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__23_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__41_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__23_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_41_ccff_tail),
		.chany_top_out(sb_1__1__21_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__21_ccff_tail));

	sb_1__1_ sb_2__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__24_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__42_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__24_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__1__22_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__22_ccff_tail));

	sb_1__1_ sb_2__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__25_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__43_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__25_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_43_ccff_tail),
		.chany_top_out(sb_1__1__23_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__23_ccff_tail));

	sb_1__1_ sb_2__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__26_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__44_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__26_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__1__24_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__24_ccff_tail));

	sb_1__1_ sb_2__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__27_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__45_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__27_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_45_ccff_tail),
		.chany_top_out(sb_1__1__25_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__25_ccff_tail));

	sb_1__1_ sb_2__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__28_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__46_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__28_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__1__26_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__26_ccff_tail));

	sb_1__1_ sb_2__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__29_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__47_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__29_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_47_ccff_tail),
		.chany_top_out(sb_1__1__27_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__27_ccff_tail));

	sb_1__1_ sb_2__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__30_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__48_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__30_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__1__28_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__28_ccff_tail));

	sb_1__1_ sb_2__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__31_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__49_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__31_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_49_ccff_tail),
		.chany_top_out(sb_1__1__29_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__29_ccff_tail));

	sb_1__1_ sb_2__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__32_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__50_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__32_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__1__30_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__30_ccff_tail));

	sb_1__1_ sb_2__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__33_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__51_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__33_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_51_ccff_tail),
		.chany_top_out(sb_1__1__31_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__31_ccff_tail));

	sb_1__1_ sb_2__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__34_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__52_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__34_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__1__32_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__32_ccff_tail));

	sb_1__1_ sb_2__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__35_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__53_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__35_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_53_ccff_tail),
		.chany_top_out(sb_1__1__33_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__33_ccff_tail));

	sb_1__1_ sb_5__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__37_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__73_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__55_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_73_ccff_tail),
		.chany_top_out(sb_1__1__34_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__34_ccff_tail));

	sb_1__1_ sb_5__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__38_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__74_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__56_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__2_ccff_tail),
		.chany_top_out(sb_1__1__35_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__35_ccff_tail));

	sb_1__1_ sb_5__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__39_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__75_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__57_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_75_ccff_tail),
		.chany_top_out(sb_1__1__36_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__36_ccff_tail));

	sb_1__1_ sb_5__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__40_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__76_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__58_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__4_ccff_tail),
		.chany_top_out(sb_1__1__37_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__37_ccff_tail));

	sb_1__1_ sb_5__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__41_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__77_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__59_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_77_ccff_tail),
		.chany_top_out(sb_1__1__38_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__38_ccff_tail));

	sb_1__1_ sb_5__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__42_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__78_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__60_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__6_ccff_tail),
		.chany_top_out(sb_1__1__39_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__39_ccff_tail));

	sb_1__1_ sb_5__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__43_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__79_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__61_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_79_ccff_tail),
		.chany_top_out(sb_1__1__40_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__40_ccff_tail));

	sb_1__1_ sb_5__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__44_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__80_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__62_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__8_ccff_tail),
		.chany_top_out(sb_1__1__41_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__41_ccff_tail));

	sb_1__1_ sb_5__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__45_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__81_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__63_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_81_ccff_tail),
		.chany_top_out(sb_1__1__42_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__42_ccff_tail));

	sb_1__1_ sb_5__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__46_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__82_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__64_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__10_ccff_tail),
		.chany_top_out(sb_1__1__43_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__43_ccff_tail));

	sb_1__1_ sb_5__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__47_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__83_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__65_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_83_ccff_tail),
		.chany_top_out(sb_1__1__44_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__44_ccff_tail));

	sb_1__1_ sb_5__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__48_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__84_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__66_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__12_ccff_tail),
		.chany_top_out(sb_1__1__45_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__45_ccff_tail));

	sb_1__1_ sb_5__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__49_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__85_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__67_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_85_ccff_tail),
		.chany_top_out(sb_1__1__46_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__46_ccff_tail));

	sb_1__1_ sb_5__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__50_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__86_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__68_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__14_ccff_tail),
		.chany_top_out(sb_1__1__47_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__47_ccff_tail));

	sb_1__1_ sb_5__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__51_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__87_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__69_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_87_ccff_tail),
		.chany_top_out(sb_1__1__48_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__48_ccff_tail));

	sb_1__1_ sb_5__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__52_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__88_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__70_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__16_ccff_tail),
		.chany_top_out(sb_1__1__49_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__49_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__49_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__49_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__49_ccff_tail));

	sb_1__1_ sb_5__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__53_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__89_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__71_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_89_ccff_tail),
		.chany_top_out(sb_1__1__50_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__50_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__50_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__50_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__50_ccff_tail));

	sb_1__1_ sb_6__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__55_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__91_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__73_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_91_ccff_tail),
		.chany_top_out(sb_1__1__51_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__51_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__51_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__51_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__51_ccff_tail));

	sb_1__1_ sb_6__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__56_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__92_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__74_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_56_ccff_tail),
		.chany_top_out(sb_1__1__52_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__52_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__52_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__52_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__52_ccff_tail));

	sb_1__1_ sb_6__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__57_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__93_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__56_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__75_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_93_ccff_tail),
		.chany_top_out(sb_1__1__53_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__53_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__53_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__53_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__53_ccff_tail));

	sb_1__1_ sb_6__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__58_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__94_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__57_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__76_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(ccff_head[4]),
		.chany_top_out(sb_1__1__54_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__54_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__54_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__54_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__54_ccff_tail));

	sb_1__1_ sb_6__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__59_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__95_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__58_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__77_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_95_ccff_tail),
		.chany_top_out(sb_1__1__55_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__55_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__55_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__55_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__55_ccff_tail));

	sb_1__1_ sb_6__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__60_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__96_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__59_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__78_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_60_ccff_tail),
		.chany_top_out(sb_1__1__56_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__56_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__56_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__56_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__56_ccff_tail));

	sb_1__1_ sb_6__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__61_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__97_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__60_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__79_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_97_ccff_tail),
		.chany_top_out(sb_1__1__57_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__57_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__57_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__57_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__57_ccff_tail));

	sb_1__1_ sb_6__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__62_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__98_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__61_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__80_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_62_ccff_tail),
		.chany_top_out(sb_1__1__58_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__58_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__58_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__58_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__58_ccff_tail));

	sb_1__1_ sb_6__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__63_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__99_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__62_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__81_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_99_ccff_tail),
		.chany_top_out(sb_1__1__59_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__59_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__59_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__59_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__59_ccff_tail));

	sb_1__1_ sb_6__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__64_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__100_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__63_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__82_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_64_ccff_tail),
		.chany_top_out(sb_1__1__60_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__60_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__60_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__60_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__60_ccff_tail));

	sb_1__1_ sb_6__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__65_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__101_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__64_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__83_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_101_ccff_tail),
		.chany_top_out(sb_1__1__61_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__61_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__61_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__61_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__61_ccff_tail));

	sb_1__1_ sb_6__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__66_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__102_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__65_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__84_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_66_ccff_tail),
		.chany_top_out(sb_1__1__62_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__62_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__62_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__62_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__62_ccff_tail));

	sb_1__1_ sb_6__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__67_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__103_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__66_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__85_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_103_ccff_tail),
		.chany_top_out(sb_1__1__63_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__63_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__63_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__63_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__63_ccff_tail));

	sb_1__1_ sb_6__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__68_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__104_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__67_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__86_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_68_ccff_tail),
		.chany_top_out(sb_1__1__64_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__64_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__64_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__64_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__64_ccff_tail));

	sb_1__1_ sb_6__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__69_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__105_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__68_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__87_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_105_ccff_tail),
		.chany_top_out(sb_1__1__65_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__65_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__65_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__65_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__65_ccff_tail));

	sb_1__1_ sb_6__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__70_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__106_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__69_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__88_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_70_ccff_tail),
		.chany_top_out(sb_1__1__66_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__66_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__66_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__66_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__66_ccff_tail));

	sb_1__1_ sb_6__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__71_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__107_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__70_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__89_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_107_ccff_tail),
		.chany_top_out(sb_1__1__67_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__67_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__67_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__67_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__67_ccff_tail));

	sb_1__1_ sb_7__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__73_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__109_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__72_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__91_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_109_ccff_tail),
		.chany_top_out(sb_1__1__68_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__68_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__68_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__68_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__68_ccff_tail));

	sb_1__1_ sb_7__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__74_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__110_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__73_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__92_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_74_ccff_tail),
		.chany_top_out(sb_1__1__69_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__69_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__69_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__69_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__69_ccff_tail));

	sb_1__1_ sb_7__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__75_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__111_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__74_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__93_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_111_ccff_tail),
		.chany_top_out(sb_1__1__70_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__70_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__70_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__70_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__70_ccff_tail));

	sb_1__1_ sb_7__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__76_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__112_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__75_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__94_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_76_ccff_tail),
		.chany_top_out(sb_1__1__71_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__71_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__71_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__71_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__71_ccff_tail));

	sb_1__1_ sb_7__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__77_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__113_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__76_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__95_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_113_ccff_tail),
		.chany_top_out(sb_1__1__72_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__72_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__72_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__72_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__72_ccff_tail));

	sb_1__1_ sb_7__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__78_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__114_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__77_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__96_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_78_ccff_tail),
		.chany_top_out(sb_1__1__73_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__73_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__73_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__73_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__73_ccff_tail));

	sb_1__1_ sb_7__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__79_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__115_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__78_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__97_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_115_ccff_tail),
		.chany_top_out(sb_1__1__74_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__74_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__74_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__74_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__74_ccff_tail));

	sb_1__1_ sb_7__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__80_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__116_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__79_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__98_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_80_ccff_tail),
		.chany_top_out(sb_1__1__75_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__75_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__75_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__75_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__75_ccff_tail));

	sb_1__1_ sb_7__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__81_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__117_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__80_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__99_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_117_ccff_tail),
		.chany_top_out(sb_1__1__76_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__76_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__76_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__76_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__76_ccff_tail));

	sb_1__1_ sb_7__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__82_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__118_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__81_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__100_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_82_ccff_tail),
		.chany_top_out(sb_1__1__77_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__77_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__77_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__77_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__77_ccff_tail));

	sb_1__1_ sb_7__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__83_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__119_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__82_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__101_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_119_ccff_tail),
		.chany_top_out(sb_1__1__78_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__78_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__78_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__78_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__78_ccff_tail));

	sb_1__1_ sb_7__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__84_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__120_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__83_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__102_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_84_ccff_tail),
		.chany_top_out(sb_1__1__79_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__79_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__79_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__79_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__79_ccff_tail));

	sb_1__1_ sb_7__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__85_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__121_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__84_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__103_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_121_ccff_tail),
		.chany_top_out(sb_1__1__80_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__80_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__80_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__80_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__80_ccff_tail));

	sb_1__1_ sb_7__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__86_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__122_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__85_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__104_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_86_ccff_tail),
		.chany_top_out(sb_1__1__81_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__81_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__81_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__81_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__81_ccff_tail));

	sb_1__1_ sb_7__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__87_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__123_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__86_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__105_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_123_ccff_tail),
		.chany_top_out(sb_1__1__82_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__82_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__82_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__82_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__82_ccff_tail));

	sb_1__1_ sb_7__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__88_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__124_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__87_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__106_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_88_ccff_tail),
		.chany_top_out(sb_1__1__83_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__83_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__83_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__83_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__83_ccff_tail));

	sb_1__1_ sb_7__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__89_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__125_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__88_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__107_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_125_ccff_tail),
		.chany_top_out(sb_1__1__84_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__84_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__84_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__84_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__84_ccff_tail));

	sb_1__1_ sb_8__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__91_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__127_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__90_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__109_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_127_ccff_tail),
		.chany_top_out(sb_1__1__85_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__85_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__85_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__85_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__85_ccff_tail));

	sb_1__1_ sb_8__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__92_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__128_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__91_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__110_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_92_ccff_tail),
		.chany_top_out(sb_1__1__86_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__86_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__86_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__86_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__86_ccff_tail));

	sb_1__1_ sb_8__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__93_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__129_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__92_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__111_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_129_ccff_tail),
		.chany_top_out(sb_1__1__87_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__87_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__87_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__87_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__87_ccff_tail));

	sb_1__1_ sb_8__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__94_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__130_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__93_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__112_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_94_ccff_tail),
		.chany_top_out(sb_1__1__88_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__88_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__88_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__88_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__88_ccff_tail));

	sb_1__1_ sb_8__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__95_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__131_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__94_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__113_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_131_ccff_tail),
		.chany_top_out(sb_1__1__89_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__89_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__89_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__89_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__89_ccff_tail));

	sb_1__1_ sb_8__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__96_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__132_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__95_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__114_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_96_ccff_tail),
		.chany_top_out(sb_1__1__90_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__90_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__90_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__90_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__90_ccff_tail));

	sb_1__1_ sb_8__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__97_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__133_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__96_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__115_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_133_ccff_tail),
		.chany_top_out(sb_1__1__91_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__91_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__91_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__91_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__91_ccff_tail));

	sb_1__1_ sb_8__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__98_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__134_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__97_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__116_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_98_ccff_tail),
		.chany_top_out(sb_1__1__92_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__92_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__92_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__92_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__92_ccff_tail));

	sb_1__1_ sb_8__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__99_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__135_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__98_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__117_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_135_ccff_tail),
		.chany_top_out(sb_1__1__93_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__93_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__93_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__93_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__93_ccff_tail));

	sb_1__1_ sb_8__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__100_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__136_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__99_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__118_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_100_ccff_tail),
		.chany_top_out(sb_1__1__94_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__94_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__94_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__94_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__94_ccff_tail));

	sb_1__1_ sb_8__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__101_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__137_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__100_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__119_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_137_ccff_tail),
		.chany_top_out(sb_1__1__95_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__95_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__95_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__95_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__95_ccff_tail));

	sb_1__1_ sb_8__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__102_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__138_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__101_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__120_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_102_ccff_tail),
		.chany_top_out(sb_1__1__96_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__96_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__96_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__96_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__96_ccff_tail));

	sb_1__1_ sb_8__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__103_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__139_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__102_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_120_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__121_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_120_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_139_ccff_tail),
		.chany_top_out(sb_1__1__97_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__97_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__97_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__97_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__97_ccff_tail));

	sb_1__1_ sb_8__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__104_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__140_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__103_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_121_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__122_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_121_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_104_ccff_tail),
		.chany_top_out(sb_1__1__98_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__98_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__98_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__98_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__98_ccff_tail));

	sb_1__1_ sb_8__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__105_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__141_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__104_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_122_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__123_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_122_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_141_ccff_tail),
		.chany_top_out(sb_1__1__99_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__99_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__99_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__99_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__99_ccff_tail));

	sb_1__1_ sb_8__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__106_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__142_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__105_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_123_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__124_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_123_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_106_ccff_tail),
		.chany_top_out(sb_1__1__100_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__100_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__100_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__100_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__100_ccff_tail));

	sb_1__1_ sb_8__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__107_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__143_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__106_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_124_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__125_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_124_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_143_ccff_tail),
		.chany_top_out(sb_1__1__101_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__101_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__101_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__101_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__101_ccff_tail));

	sb_1__1_ sb_9__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__109_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__145_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__108_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_126_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__127_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_126_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_145_ccff_tail),
		.chany_top_out(sb_1__1__102_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__102_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__102_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__102_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__102_ccff_tail));

	sb_1__1_ sb_9__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__110_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__146_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__109_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_127_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__128_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_127_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_110_ccff_tail),
		.chany_top_out(sb_1__1__103_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__103_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__103_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__103_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__103_ccff_tail));

	sb_1__1_ sb_9__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__111_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__147_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__110_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_128_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__129_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_128_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_147_ccff_tail),
		.chany_top_out(sb_1__1__104_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__104_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__104_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__104_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__104_ccff_tail));

	sb_1__1_ sb_9__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__112_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__148_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__111_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_129_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__130_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_129_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_112_ccff_tail),
		.chany_top_out(sb_1__1__105_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__105_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__105_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__105_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__105_ccff_tail));

	sb_1__1_ sb_9__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__113_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__149_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__112_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_130_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__131_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_130_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_149_ccff_tail),
		.chany_top_out(sb_1__1__106_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__106_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__106_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__106_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__106_ccff_tail));

	sb_1__1_ sb_9__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__114_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__150_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__113_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_131_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__132_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_131_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_114_ccff_tail),
		.chany_top_out(sb_1__1__107_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__107_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__107_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__107_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__107_ccff_tail));

	sb_1__1_ sb_9__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__115_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__151_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__114_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_132_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__133_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_132_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_151_ccff_tail),
		.chany_top_out(sb_1__1__108_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__108_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__108_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__108_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__108_ccff_tail));

	sb_1__1_ sb_9__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__116_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__152_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__115_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_133_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__134_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_133_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_116_ccff_tail),
		.chany_top_out(sb_1__1__109_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__109_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__109_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__109_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__109_ccff_tail));

	sb_1__1_ sb_9__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__117_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__153_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__116_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_134_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__135_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_134_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_153_ccff_tail),
		.chany_top_out(sb_1__1__110_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__110_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__110_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__110_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__110_ccff_tail));

	sb_1__1_ sb_9__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__118_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__154_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__117_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_135_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__136_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_135_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_118_ccff_tail),
		.chany_top_out(sb_1__1__111_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__111_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__111_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__111_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__111_ccff_tail));

	sb_1__1_ sb_9__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__119_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__155_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__118_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_136_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__137_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_136_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_155_ccff_tail),
		.chany_top_out(sb_1__1__112_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__112_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__112_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__112_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__112_ccff_tail));

	sb_1__1_ sb_9__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__120_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__156_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__119_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_137_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__138_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_137_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_120_ccff_tail),
		.chany_top_out(sb_1__1__113_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__113_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__113_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__113_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__113_ccff_tail));

	sb_1__1_ sb_9__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__121_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__157_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__120_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_138_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__139_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_138_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_157_ccff_tail),
		.chany_top_out(sb_1__1__114_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__114_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__114_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__114_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__114_ccff_tail));

	sb_1__1_ sb_9__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__122_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__158_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__121_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_139_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__140_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_139_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_122_ccff_tail),
		.chany_top_out(sb_1__1__115_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__115_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__115_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__115_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__115_ccff_tail));

	sb_1__1_ sb_9__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__123_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__159_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__122_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_140_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__141_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_140_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_159_ccff_tail),
		.chany_top_out(sb_1__1__116_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__116_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__116_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__116_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__116_ccff_tail));

	sb_1__1_ sb_9__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__124_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__160_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__123_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_141_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__142_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_141_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_124_ccff_tail),
		.chany_top_out(sb_1__1__117_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__117_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__117_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__117_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__117_ccff_tail));

	sb_1__1_ sb_9__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__125_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__161_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__124_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_142_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__143_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_142_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_161_ccff_tail),
		.chany_top_out(sb_1__1__118_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__118_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__118_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__118_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__118_ccff_tail));

	sb_1__1_ sb_12__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__127_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__181_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__126_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_162_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__163_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_181_ccff_tail),
		.chany_top_out(sb_1__1__119_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__119_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__119_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__119_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__119_ccff_tail));

	sb_1__1_ sb_12__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__128_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__182_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__127_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_163_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__164_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__20_ccff_tail),
		.chany_top_out(sb_1__1__120_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__120_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__120_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__120_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__120_ccff_tail));

	sb_1__1_ sb_12__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__129_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__183_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__128_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_164_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__165_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_183_ccff_tail),
		.chany_top_out(sb_1__1__121_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__121_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__121_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__121_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__121_ccff_tail));

	sb_1__1_ sb_12__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__130_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__184_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__129_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_165_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__166_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__22_ccff_tail),
		.chany_top_out(sb_1__1__122_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__122_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__122_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__122_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__122_ccff_tail));

	sb_1__1_ sb_12__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__131_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__185_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__130_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_166_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__167_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_185_ccff_tail),
		.chany_top_out(sb_1__1__123_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__123_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__123_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__123_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__123_ccff_tail));

	sb_1__1_ sb_12__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__132_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__186_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__131_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_167_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__168_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__24_ccff_tail),
		.chany_top_out(sb_1__1__124_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__124_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__124_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__124_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__124_ccff_tail));

	sb_1__1_ sb_12__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__133_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__187_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__132_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_168_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__169_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_187_ccff_tail),
		.chany_top_out(sb_1__1__125_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__125_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__125_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__125_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__125_ccff_tail));

	sb_1__1_ sb_12__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__134_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__188_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__133_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_169_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__170_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__26_ccff_tail),
		.chany_top_out(sb_1__1__126_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__126_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__126_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__126_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__126_ccff_tail));

	sb_1__1_ sb_12__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__135_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__189_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__134_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_170_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__171_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_189_ccff_tail),
		.chany_top_out(sb_1__1__127_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__127_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__127_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__127_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__127_ccff_tail));

	sb_1__1_ sb_12__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__136_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__190_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__135_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_171_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__172_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__28_ccff_tail),
		.chany_top_out(sb_1__1__128_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__128_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__128_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__128_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__128_ccff_tail));

	sb_1__1_ sb_12__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__137_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__191_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__136_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_172_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__173_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_191_ccff_tail),
		.chany_top_out(sb_1__1__129_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__129_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__129_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__129_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__129_ccff_tail));

	sb_1__1_ sb_12__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__138_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__192_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__137_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_173_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__174_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(ccff_head[9]),
		.chany_top_out(sb_1__1__130_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__130_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__130_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__130_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__130_ccff_tail));

	sb_1__1_ sb_12__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__139_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__193_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__138_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_174_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__175_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_193_ccff_tail),
		.chany_top_out(sb_1__1__131_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__131_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__131_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__131_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__131_ccff_tail));

	sb_1__1_ sb_12__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__140_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__194_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__139_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_175_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__176_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__32_ccff_tail),
		.chany_top_out(sb_1__1__132_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__132_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__132_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__132_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__132_ccff_tail));

	sb_1__1_ sb_12__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__141_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__195_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__140_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_176_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__177_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_195_ccff_tail),
		.chany_top_out(sb_1__1__133_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__133_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__133_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__133_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__133_ccff_tail));

	sb_1__1_ sb_12__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__142_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__196_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__141_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_177_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__178_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__34_ccff_tail),
		.chany_top_out(sb_1__1__134_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__134_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__134_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__134_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__134_ccff_tail));

	sb_1__1_ sb_12__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__143_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__197_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__142_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_178_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__179_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_197_ccff_tail),
		.chany_top_out(sb_1__1__135_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__135_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__135_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__135_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__135_ccff_tail));

	sb_1__1_ sb_13__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__145_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__199_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__144_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_180_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__181_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_180_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_199_ccff_tail),
		.chany_top_out(sb_1__1__136_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__136_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__136_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__136_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__136_ccff_tail));

	sb_1__1_ sb_13__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__146_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__200_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__145_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_181_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__182_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_181_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_164_ccff_tail),
		.chany_top_out(sb_1__1__137_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__137_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__137_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__137_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__137_ccff_tail));

	sb_1__1_ sb_13__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__147_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__201_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__146_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_182_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__183_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_182_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_201_ccff_tail),
		.chany_top_out(sb_1__1__138_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__138_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__138_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__138_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__138_ccff_tail));

	sb_1__1_ sb_13__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__148_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__202_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__147_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_183_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__184_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_183_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_166_ccff_tail),
		.chany_top_out(sb_1__1__139_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__139_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__139_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__139_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__139_ccff_tail));

	sb_1__1_ sb_13__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__149_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__203_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__148_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_184_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__185_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_184_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_203_ccff_tail),
		.chany_top_out(sb_1__1__140_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__140_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__140_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__140_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__140_ccff_tail));

	sb_1__1_ sb_13__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__150_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__204_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__149_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_185_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__186_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_185_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_168_ccff_tail),
		.chany_top_out(sb_1__1__141_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__141_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__141_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__141_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__141_ccff_tail));

	sb_1__1_ sb_13__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__151_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__205_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__150_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_186_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__187_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_186_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_205_ccff_tail),
		.chany_top_out(sb_1__1__142_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__142_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__142_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__142_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__142_ccff_tail));

	sb_1__1_ sb_13__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__152_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__206_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__151_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_187_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__188_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_187_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_170_ccff_tail),
		.chany_top_out(sb_1__1__143_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__143_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__143_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__143_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__143_ccff_tail));

	sb_1__1_ sb_13__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__153_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__207_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__152_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_188_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__189_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_188_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_207_ccff_tail),
		.chany_top_out(sb_1__1__144_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__144_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__144_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__144_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__144_ccff_tail));

	sb_1__1_ sb_13__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__154_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__208_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__153_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_189_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__190_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_189_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_172_ccff_tail),
		.chany_top_out(sb_1__1__145_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__145_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__145_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__145_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__145_ccff_tail));

	sb_1__1_ sb_13__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__155_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__209_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__154_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_190_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__191_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_190_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_209_ccff_tail),
		.chany_top_out(sb_1__1__146_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__146_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__146_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__146_chanx_left_out[0:63]),
		.ccff_tail(ccff_tail[7]));

	sb_1__1_ sb_13__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__156_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__210_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__155_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_191_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__192_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_191_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_174_ccff_tail),
		.chany_top_out(sb_1__1__147_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__147_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__147_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__147_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__147_ccff_tail));

	sb_1__1_ sb_13__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__157_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__211_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__156_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_192_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__193_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_192_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_211_ccff_tail),
		.chany_top_out(sb_1__1__148_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__148_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__148_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__148_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__148_ccff_tail));

	sb_1__1_ sb_13__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__158_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__212_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__157_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_193_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__194_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_193_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_176_ccff_tail),
		.chany_top_out(sb_1__1__149_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__149_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__149_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__149_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__149_ccff_tail));

	sb_1__1_ sb_13__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__159_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__213_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__158_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_194_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__195_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_194_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_213_ccff_tail),
		.chany_top_out(sb_1__1__150_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__150_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__150_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__150_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__150_ccff_tail));

	sb_1__1_ sb_13__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__160_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__214_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__159_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_195_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__196_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_195_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_178_ccff_tail),
		.chany_top_out(sb_1__1__151_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__151_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__151_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__151_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__151_ccff_tail));

	sb_1__1_ sb_13__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__161_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.chanx_right_in(cbx_1__0__215_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__160_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_196_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__197_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_196_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_215_ccff_tail),
		.chany_top_out(sb_1__1__152_chany_top_out[0:63]),
		.chanx_right_out(sb_1__1__152_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__1__152_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__1__152_chanx_left_out[0:63]),
		.ccff_tail(sb_1__1__152_ccff_tail));

	sb_1__18_ sb_1__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__1_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__0_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_1_ccff_tail),
		.chanx_right_out(sb_1__18__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__0_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__0_ccff_tail));

	sb_1__18_ sb_2__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__2_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__1_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_2_ccff_tail),
		.chanx_right_out(sb_1__18__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__1_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__1_ccff_tail));

	sb_1__18_ sb_5__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__4_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__3_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_5_ccff_tail),
		.chanx_right_out(sb_1__18__2_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__2_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__2_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__2_ccff_tail));

	sb_1__18_ sb_6__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__5_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__71_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__4_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_6_ccff_tail),
		.chanx_right_out(sb_1__18__3_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__3_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__3_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__3_ccff_tail));

	sb_1__18_ sb_7__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__6_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__89_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__5_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_7_ccff_tail),
		.chanx_right_out(sb_1__18__4_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__4_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__4_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__4_ccff_tail));

	sb_1__18_ sb_8__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__7_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__107_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_125_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__6_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_125_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_8_ccff_tail),
		.chanx_right_out(sb_1__18__5_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__5_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__5_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__5_ccff_tail));

	sb_1__18_ sb_9__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__8_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__125_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_143_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__7_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_143_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_9_ccff_tail),
		.chanx_right_out(sb_1__18__6_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__6_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__6_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__6_ccff_tail));

	sb_1__18_ sb_12__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__10_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__143_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_179_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__9_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_12_ccff_tail),
		.chanx_right_out(sb_1__18__7_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__7_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__7_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__7_ccff_tail));

	sb_1__18_ sb_13__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__11_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_1__1__161_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_197_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__10_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_197_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_13_ccff_tail),
		.chanx_right_out(sb_1__18__8_chanx_right_out[0:63]),
		.chany_bottom_out(sb_1__18__8_chany_bottom_out[0:63]),
		.chanx_left_out(sb_1__18__8_chanx_left_out[0:63]),
		.ccff_tail(sb_1__18__8_ccff_tail));

	sb_3__0_ sb_3__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__0__0_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__36_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_3__0__0_chany_top_out[0:63]),
		.chanx_right_out(sb_3__0__0_chanx_right_out[0:63]),
		.chanx_left_out(sb_3__0__0_chanx_left_out[0:63]),
		.ccff_tail(sb_3__0__0_ccff_tail));

	sb_3__0_ sb_10__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__0__1_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__144_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_126_ccff_tail),
		.chany_top_out(sb_3__0__1_chany_top_out[0:63]),
		.chanx_right_out(sb_3__0__1_chanx_right_out[0:63]),
		.chanx_left_out(sb_3__0__1_chanx_left_out[0:63]),
		.ccff_tail(sb_3__0__1_ccff_tail));

	sb_3__1_ sb_3__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__0_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__0_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__37_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__1_ccff_tail),
		.chany_top_out(sb_3__1__0_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__0_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__0_ccff_tail));

	sb_3__1_ sb_3__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__0_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__0_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__38_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_3__1__1_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__1_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__1_ccff_tail));

	sb_3__1_ sb_3__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__1_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__1_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_1_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__39_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__3_ccff_tail),
		.chany_top_out(sb_3__1__2_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__2_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__2_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__2_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__2_ccff_tail));

	sb_3__1_ sb_3__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__1_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__1_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_1_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__40_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_3__1__3_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__3_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__3_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__3_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__3_ccff_tail));

	sb_3__1_ sb_3__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__2_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__2_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_2_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__41_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__5_ccff_tail),
		.chany_top_out(sb_3__1__4_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__4_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__4_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__4_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__4_ccff_tail));

	sb_3__1_ sb_3__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__2_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__2_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_2_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__42_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_24_ccff_tail),
		.chany_top_out(sb_3__1__5_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__5_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__5_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__5_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__5_ccff_tail));

	sb_3__1_ sb_3__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__3_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__3_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_3_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__43_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__7_ccff_tail),
		.chany_top_out(sb_3__1__6_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__6_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__6_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__6_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__6_ccff_tail));

	sb_3__1_ sb_3__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__3_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__3_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_3_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__44_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_26_ccff_tail),
		.chany_top_out(sb_3__1__7_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__7_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__7_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__7_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__7_ccff_tail));

	sb_3__1_ sb_3__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__4_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__4_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_4_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__45_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__9_ccff_tail),
		.chany_top_out(sb_3__1__8_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__8_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__8_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__8_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__8_ccff_tail));

	sb_3__1_ sb_3__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__4_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__4_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_4_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__46_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_28_ccff_tail),
		.chany_top_out(sb_3__1__9_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__9_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__9_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__9_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__9_ccff_tail));

	sb_3__1_ sb_3__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__5_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__5_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_5_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__47_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__11_ccff_tail),
		.chany_top_out(sb_3__1__10_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__10_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__10_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__10_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__10_ccff_tail));

	sb_3__1_ sb_3__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__5_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__5_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_5_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__48_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_30_ccff_tail),
		.chany_top_out(sb_3__1__11_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__11_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__11_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__11_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__11_ccff_tail));

	sb_3__1_ sb_3__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__6_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__6_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_6_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__49_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__13_ccff_tail),
		.chany_top_out(sb_3__1__12_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__12_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__12_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__12_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__12_ccff_tail));

	sb_3__1_ sb_3__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__6_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__6_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_6_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__50_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_32_ccff_tail),
		.chany_top_out(sb_3__1__13_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__13_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__13_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__13_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__13_ccff_tail));

	sb_3__1_ sb_3__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__7_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__7_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_7_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__51_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__15_ccff_tail),
		.chany_top_out(sb_3__1__14_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__14_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__14_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__14_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__14_ccff_tail));

	sb_3__1_ sb_3__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__7_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__7_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_7_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__52_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(ccff_head[11]),
		.chany_top_out(sb_3__1__15_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__15_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__15_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__15_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__15_ccff_tail));

	sb_3__1_ sb_3__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__8_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__8_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_8_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__53_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__17_ccff_tail),
		.chany_top_out(sb_3__1__16_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__16_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__16_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__16_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__16_ccff_tail));

	sb_3__1_ sb_10__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__9_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__9_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_9_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_144_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__145_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_144_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__19_ccff_tail),
		.chany_top_out(sb_3__1__17_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__17_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__17_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__17_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__17_ccff_tail));

	sb_3__1_ sb_10__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__8_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__9_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_9_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_145_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__146_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_145_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_128_ccff_tail),
		.chany_top_out(sb_3__1__18_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__18_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__18_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__18_chanx_left_out[0:63]),
		.ccff_tail(ccff_tail[2]));

	sb_3__1_ sb_10__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__10_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__10_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_10_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_146_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__147_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_146_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__21_ccff_tail),
		.chany_top_out(sb_3__1__19_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__19_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__19_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__19_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__19_ccff_tail));

	sb_3__1_ sb_10__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__9_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__10_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_10_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_147_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__148_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_147_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_130_ccff_tail),
		.chany_top_out(sb_3__1__20_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__20_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__20_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__20_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__20_ccff_tail));

	sb_3__1_ sb_10__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__11_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__11_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_11_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_148_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__149_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_148_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__23_ccff_tail),
		.chany_top_out(sb_3__1__21_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__21_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__21_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__21_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__21_ccff_tail));

	sb_3__1_ sb_10__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__10_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__11_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_11_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_149_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__150_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_149_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_132_ccff_tail),
		.chany_top_out(sb_3__1__22_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__22_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__22_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__22_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__22_ccff_tail));

	sb_3__1_ sb_10__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__12_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__12_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_12_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_150_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__151_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_150_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__25_ccff_tail),
		.chany_top_out(sb_3__1__23_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__23_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__23_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__23_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__23_ccff_tail));

	sb_3__1_ sb_10__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__11_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__12_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_12_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_151_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__152_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_151_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_134_ccff_tail),
		.chany_top_out(sb_3__1__24_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__24_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__24_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__24_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__24_ccff_tail));

	sb_3__1_ sb_10__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__13_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__13_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_13_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_152_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__153_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_152_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__27_ccff_tail),
		.chany_top_out(sb_3__1__25_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__25_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__25_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__25_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__25_ccff_tail));

	sb_3__1_ sb_10__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__12_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__13_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_13_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_153_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__154_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_153_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_136_ccff_tail),
		.chany_top_out(sb_3__1__26_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__26_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__26_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__26_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__26_ccff_tail));

	sb_3__1_ sb_10__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__14_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__14_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_14_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_154_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__155_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_154_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__29_ccff_tail),
		.chany_top_out(sb_3__1__27_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__27_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__27_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__27_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__27_ccff_tail));

	sb_3__1_ sb_10__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__13_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__14_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_14_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_155_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__156_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_155_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_138_ccff_tail),
		.chany_top_out(sb_3__1__28_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__28_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__28_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__28_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__28_ccff_tail));

	sb_3__1_ sb_10__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__15_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__15_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_15_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_156_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__157_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_156_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__31_ccff_tail),
		.chany_top_out(sb_3__1__29_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__29_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__29_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__29_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__29_ccff_tail));

	sb_3__1_ sb_10__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__14_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__15_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_15_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_157_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__158_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_157_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_140_ccff_tail),
		.chany_top_out(sb_3__1__30_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__30_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__30_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__30_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__30_ccff_tail));

	sb_3__1_ sb_10__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__16_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__16_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_16_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_158_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__159_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_158_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__33_ccff_tail),
		.chany_top_out(sb_3__1__31_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__31_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__31_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__31_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__31_ccff_tail));

	sb_3__1_ sb_10__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__1__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_lower),
		.chanx_right_in(cbx_4__2__15_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__16_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_16_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_159_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__160_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_159_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_142_ccff_tail),
		.chany_top_out(sb_3__1__32_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__32_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__32_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__32_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__32_ccff_tail));

	sb_3__1_ sb_10__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_lower),
		.chanx_right_in(cbx_4__1__17_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_upper),
		.chany_bottom_in(cby_3__1__17_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_17_left_width_0_height_0_subtile_0__pin_data_out_2_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_160_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__161_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_160_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(cby_4__1__35_ccff_tail),
		.chany_top_out(sb_3__1__33_chany_top_out[0:63]),
		.chanx_right_out(sb_3__1__33_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__1__33_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__1__33_chanx_left_out[0:63]),
		.ccff_tail(sb_3__1__33_ccff_tail));

	sb_3__18_ sb_3__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_4__18__0_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_1_subtile_0__pin_data_out_5_(grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__8_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_8_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__2_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_3_ccff_tail),
		.chanx_right_out(sb_3__18__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__18__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__18__0_chanx_left_out[0:63]),
		.ccff_tail(sb_3__18__0_ccff_tail));

	sb_3__18_ sb_10__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_4__18__1_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_1_subtile_0__pin_data_out_5_(grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_upper),
		.chany_bottom_in(cby_3__2__17_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_1_subtile_0__pin_data_out_3_(grid_memory_17_left_width_0_height_1_subtile_0__pin_data_out_3_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_161_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__8_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_161_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_top_top_10_ccff_tail),
		.chanx_right_out(sb_3__18__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_3__18__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_3__18__1_chanx_left_out[0:63]),
		.ccff_tail(sb_3__18__1_ccff_tail));

	sb_4__0_ sb_4__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__54_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_4__0__0_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_36_ccff_tail),
		.chany_top_out(sb_4__0__0_chany_top_out[0:63]),
		.chanx_right_out(sb_4__0__0_chanx_right_out[0:63]),
		.chanx_left_out(sb_4__0__0_chanx_left_out[0:63]),
		.ccff_tail(sb_4__0__0_ccff_tail));

	sb_4__0_ sb_11__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__18_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__162_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_4__0__1_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_9_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_144_ccff_tail),
		.chany_top_out(sb_4__0__1_chany_top_out[0:63]),
		.chanx_right_out(sb_4__0__1_chanx_right_out[0:63]),
		.chanx_left_out(sb_4__0__1_chanx_left_out[0:63]),
		.ccff_tail(sb_4__0__1_ccff_tail));

	sb_4__1_ sb_4__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__55_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__0_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__0_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_0_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_55_ccff_tail),
		.chany_top_out(sb_4__1__0_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__0_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__0_ccff_tail));

	sb_4__1_ sb_4__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__56_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__1_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__0_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_1_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_38_ccff_tail),
		.chany_top_out(sb_4__1__1_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__1_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__1_ccff_tail));

	sb_4__1_ sb_4__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__57_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__2_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_1_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__1_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_1_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_1_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_57_ccff_tail),
		.chany_top_out(sb_4__1__2_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__2_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__2_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__2_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__2_ccff_tail));

	sb_4__1_ sb_4__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__58_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__3_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_1_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__1_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_2_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_1_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_40_ccff_tail),
		.chany_top_out(sb_4__1__3_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__3_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__3_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__3_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__3_ccff_tail));

	sb_4__1_ sb_4__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__59_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__4_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_2_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__2_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_2_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_59_ccff_tail),
		.chany_top_out(sb_4__1__4_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__4_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__4_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__4_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__4_ccff_tail));

	sb_4__1_ sb_4__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__60_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__5_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_2_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__2_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_3_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_2_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_42_ccff_tail),
		.chany_top_out(sb_4__1__5_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__5_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__5_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__5_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__5_ccff_tail));

	sb_4__1_ sb_4__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__61_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__6_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_3_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__3_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_3_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_3_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(ccff_head[6]),
		.chany_top_out(sb_4__1__6_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__6_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__6_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__6_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__6_ccff_tail));

	sb_4__1_ sb_4__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__62_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__7_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_3_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__3_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_4_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_3_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_44_ccff_tail),
		.chany_top_out(sb_4__1__7_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__7_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__7_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__7_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__7_ccff_tail));

	sb_4__1_ sb_4__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__63_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__8_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_4_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__4_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_4_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_4_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_63_ccff_tail),
		.chany_top_out(sb_4__1__8_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__8_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__8_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__8_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__8_ccff_tail));

	sb_4__1_ sb_4__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__64_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__9_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_4_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__4_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_5_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_4_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_46_ccff_tail),
		.chany_top_out(sb_4__1__9_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__9_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__9_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__9_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__9_ccff_tail));

	sb_4__1_ sb_4__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__65_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__10_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_5_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__5_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_5_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_5_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_65_ccff_tail),
		.chany_top_out(sb_4__1__10_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__10_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__10_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__10_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__10_ccff_tail));

	sb_4__1_ sb_4__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__66_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__11_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_5_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__5_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_6_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_5_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_48_ccff_tail),
		.chany_top_out(sb_4__1__11_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__11_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__11_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__11_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__11_ccff_tail));

	sb_4__1_ sb_4__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__67_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__12_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_6_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__6_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_6_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_6_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_67_ccff_tail),
		.chany_top_out(sb_4__1__12_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__12_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__12_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__12_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__12_ccff_tail));

	sb_4__1_ sb_4__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__68_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__13_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_6_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__6_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_7_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_6_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_50_ccff_tail),
		.chany_top_out(sb_4__1__13_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__13_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__13_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__13_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__13_ccff_tail));

	sb_4__1_ sb_4__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__69_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__14_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_7_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__7_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_7_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_7_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_69_ccff_tail),
		.chany_top_out(sb_4__1__14_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__14_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__14_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__14_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__14_ccff_tail));

	sb_4__1_ sb_4__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__70_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__15_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_7_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__7_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_8_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_7_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_52_ccff_tail),
		.chany_top_out(sb_4__1__15_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__15_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__15_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__15_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__15_ccff_tail));

	sb_4__1_ sb_4__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__71_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__16_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_8_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__8_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_8_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_8_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_71_ccff_tail),
		.chany_top_out(sb_4__1__16_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__16_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__16_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__16_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__16_ccff_tail));

	sb_4__1_ sb_11__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__19_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__163_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_162_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__18_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_9_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__9_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_9_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_9_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_163_ccff_tail),
		.chany_top_out(sb_4__1__17_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__17_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__17_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__17_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__17_ccff_tail));

	sb_4__1_ sb_11__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__20_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__164_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_163_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__19_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_9_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__8_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_10_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_9_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_146_ccff_tail),
		.chany_top_out(sb_4__1__18_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__18_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__18_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__18_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__18_ccff_tail));

	sb_4__1_ sb_11__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__21_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__165_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_164_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__20_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_10_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__10_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_10_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_10_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_165_ccff_tail),
		.chany_top_out(sb_4__1__19_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__19_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__19_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__19_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__19_ccff_tail));

	sb_4__1_ sb_11__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__22_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__166_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_165_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__21_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_10_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__9_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_11_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_10_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_148_ccff_tail),
		.chany_top_out(sb_4__1__20_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__20_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__20_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__20_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__20_ccff_tail));

	sb_4__1_ sb_11__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__23_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__167_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_166_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__22_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_11_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__11_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_11_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_11_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_167_ccff_tail),
		.chany_top_out(sb_4__1__21_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__21_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__21_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__21_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__21_ccff_tail));

	sb_4__1_ sb_11__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__24_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__168_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_167_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__23_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_11_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__10_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_12_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_11_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_150_ccff_tail),
		.chany_top_out(sb_4__1__22_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__22_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__22_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__22_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__22_ccff_tail));

	sb_4__1_ sb_11__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__25_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__169_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_168_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__24_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_12_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__12_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_12_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_12_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_169_ccff_tail),
		.chany_top_out(sb_4__1__23_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__23_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__23_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__23_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__23_ccff_tail));

	sb_4__1_ sb_11__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__26_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__170_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_169_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__25_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_12_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__11_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_13_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_12_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_152_ccff_tail),
		.chany_top_out(sb_4__1__24_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__24_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__24_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__24_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__24_ccff_tail));

	sb_4__1_ sb_11__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__27_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__171_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_170_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__26_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_13_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__13_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_13_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_13_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_171_ccff_tail),
		.chany_top_out(sb_4__1__25_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__25_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__25_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__25_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__25_ccff_tail));

	sb_4__1_ sb_11__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__28_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__172_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_171_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__27_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_13_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__12_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_14_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_13_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_154_ccff_tail),
		.chany_top_out(sb_4__1__26_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__26_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__26_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__26_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__26_ccff_tail));

	sb_4__1_ sb_11__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__29_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__173_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_172_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__28_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_14_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__14_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_14_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_14_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_173_ccff_tail),
		.chany_top_out(sb_4__1__27_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__27_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__27_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__27_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__27_ccff_tail));

	sb_4__1_ sb_11__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__30_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__174_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_173_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__29_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_14_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__13_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_15_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_14_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_156_ccff_tail),
		.chany_top_out(sb_4__1__28_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__28_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__28_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__28_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__28_ccff_tail));

	sb_4__1_ sb_11__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__31_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__175_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_174_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__30_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_15_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__15_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_15_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_15_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_175_ccff_tail),
		.chany_top_out(sb_4__1__29_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__29_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__29_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__29_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__29_ccff_tail));

	sb_4__1_ sb_11__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__32_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__176_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_175_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__31_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_15_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__14_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_16_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_15_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_158_ccff_tail),
		.chany_top_out(sb_4__1__30_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__30_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__30_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__30_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__30_ccff_tail));

	sb_4__1_ sb_11__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__33_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__177_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_176_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__32_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_16_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__16_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_16_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_16_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_177_ccff_tail),
		.chany_top_out(sb_4__1__31_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__31_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__31_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__31_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__31_ccff_tail));

	sb_4__1_ sb_11__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__34_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_lower),
		.chanx_right_in(cbx_1__0__178_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_177_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__33_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_16_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__2__15_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_17_bottom_width_0_height_0_subtile_0__pin_data_out_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_16_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_clb_160_ccff_tail),
		.chany_top_out(sb_4__1__32_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__32_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__32_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__32_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__32_ccff_tail));

	sb_4__1_ sb_11__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__35_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_lower),
		.chanx_right_in(cbx_1__0__179_chanx_left_out[0:63]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_178_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__34_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_17_right_width_0_height_0_subtile_0__pin_data_out_6_upper),
		.chanx_left_in(cbx_4__1__17_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_1_subtile_0__pin_data_out_1_(grid_memory_17_bottom_width_0_height_1_subtile_0__pin_data_out_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_17_top_width_0_height_0_subtile_0__pin_data_out_4_lower),
		.ccff_head(grid_clb_179_ccff_tail),
		.chany_top_out(sb_4__1__33_chany_top_out[0:63]),
		.chanx_right_out(sb_4__1__33_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__1__33_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__1__33_chanx_left_out[0:63]),
		.ccff_tail(sb_4__1__33_ccff_tail));

	sb_4__18_ sb_4__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__3_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__17_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_8_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__18__0_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_1_subtile_0__pin_data_out_5_(grid_memory_8_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_io_top_top_4_ccff_tail),
		.chanx_right_out(sb_4__18__0_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__18__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__18__0_chanx_left_out[0:63]),
		.ccff_tail(sb_4__18__0_ccff_tail));

	sb_4__18_ sb_11__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__18__9_chanx_left_out[0:63]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_179_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.chany_bottom_in(cby_4__1__35_chany_top_out[0:63]),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_data_out_7_(grid_memory_17_right_width_0_height_1_subtile_0__pin_data_out_7_upper),
		.chanx_left_in(cbx_4__18__1_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_1_subtile_0__pin_data_out_5_(grid_memory_17_top_width_0_height_1_subtile_0__pin_data_out_5_lower),
		.ccff_head(grid_io_top_top_11_ccff_tail),
		.chanx_right_out(sb_4__18__1_chanx_right_out[0:63]),
		.chany_bottom_out(sb_4__18__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_4__18__1_chanx_left_out[0:63]),
		.ccff_tail(sb_4__18__1_ccff_tail));

	sb_14__0_ sb_14__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__0_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_left_in(cbx_1__0__198_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_clb_180_ccff_tail),
		.chany_top_out(sb_14__0__0_chany_top_out[0:63]),
		.chanx_left_out(sb_14__0__0_chanx_left_out[0:63]),
		.ccff_tail(sb_14__0__0_ccff_tail));

	sb_14__1_ sb_14__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__1_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__0_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_198_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__199_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_198_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_198_ccff_tail),
		.chany_top_out(sb_14__1__0_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__0_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__0_ccff_tail));

	sb_14__1_ sb_14__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__2_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__1_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_199_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__200_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_199_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_182_ccff_tail),
		.chany_top_out(sb_14__1__1_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__1_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__1_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__1_ccff_tail));

	sb_14__1_ sb_14__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__3_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__2_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_200_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__201_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_200_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_200_ccff_tail),
		.chany_top_out(sb_14__1__2_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__2_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__2_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__2_ccff_tail));

	sb_14__1_ sb_14__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__4_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__3_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_201_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__202_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_201_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_184_ccff_tail),
		.chany_top_out(sb_14__1__3_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__3_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__3_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__3_ccff_tail));

	sb_14__1_ sb_14__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__5_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__4_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_202_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__203_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_202_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_202_ccff_tail),
		.chany_top_out(sb_14__1__4_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__4_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__4_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__4_ccff_tail));

	sb_14__1_ sb_14__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__6_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__5_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_203_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__204_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_203_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_186_ccff_tail),
		.chany_top_out(sb_14__1__5_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__5_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__5_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__5_ccff_tail));

	sb_14__1_ sb_14__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__7_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__6_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_204_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__205_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_204_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_204_ccff_tail),
		.chany_top_out(sb_14__1__6_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__6_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__6_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__6_ccff_tail));

	sb_14__1_ sb_14__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__8_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__7_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_205_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__206_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_205_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_188_ccff_tail),
		.chany_top_out(sb_14__1__7_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__7_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__7_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__7_ccff_tail));

	sb_14__1_ sb_14__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__9_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__8_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_206_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__207_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_206_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_206_ccff_tail),
		.chany_top_out(sb_14__1__8_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__8_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__8_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__8_ccff_tail));

	sb_14__1_ sb_14__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__10_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__9_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_207_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__208_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_207_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_190_ccff_tail),
		.chany_top_out(sb_14__1__9_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__9_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__9_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__9_ccff_tail));

	sb_14__1_ sb_14__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__11_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__10_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_208_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__209_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_208_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_208_ccff_tail),
		.chany_top_out(sb_14__1__10_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__10_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__10_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__10_ccff_tail));

	sb_14__1_ sb_14__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__12_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__11_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_209_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__210_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_209_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_192_ccff_tail),
		.chany_top_out(sb_14__1__11_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__11_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__11_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__11_ccff_tail));

	sb_14__1_ sb_14__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__13_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__12_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_210_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__211_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_210_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_210_ccff_tail),
		.chany_top_out(sb_14__1__12_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__12_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__12_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__12_ccff_tail));

	sb_14__1_ sb_14__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__14_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__13_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_211_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__212_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_211_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_194_ccff_tail),
		.chany_top_out(sb_14__1__13_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__13_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__13_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__13_ccff_tail));

	sb_14__1_ sb_14__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__15_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__14_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_212_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__213_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_212_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_212_ccff_tail),
		.chany_top_out(sb_14__1__14_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__14_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__14_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__14_ccff_tail));

	sb_14__1_ sb_14__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__16_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__15_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_213_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__214_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_213_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_196_ccff_tail),
		.chany_top_out(sb_14__1__15_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__15_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__15_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__15_ccff_tail));

	sb_14__1_ sb_14__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_14__1__17_chany_bottom_out[0:63]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_14__1__16_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_214_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__0__215_chanx_right_out[0:63]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_214_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_clb_214_ccff_tail),
		.chany_top_out(sb_14__1__16_chany_top_out[0:63]),
		.chany_bottom_out(sb_14__1__16_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__1__16_chanx_left_out[0:63]),
		.ccff_tail(sb_14__1__16_ccff_tail));

	sb_14__18_ sb_14__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_14__1__17_chany_top_out[0:63]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_4_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_5_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_6_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_215_right_width_0_height_0_subtile_0__pin_O_7_upper),
		.chanx_left_in(cbx_1__18__11_chanx_right_out[0:63]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_215_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.ccff_head(grid_io_right_right_0_ccff_tail),
		.chany_bottom_out(sb_14__18__0_chany_bottom_out[0:63]),
		.chanx_left_out(sb_14__18__0_chanx_left_out[0:63]),
		.ccff_tail(sb_14__18__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_1__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_1__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_1__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_1__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_1__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__0_ cbx_1__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(ccff_tail[4]));

	cbx_1__0_ cbx_1__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__7_ccff_tail));

	cbx_1__0_ cbx_1__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__0__8_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__8_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__8_ccff_tail));

	cbx_1__0_ cbx_1__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__0__9_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__9_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__9_ccff_tail));

	cbx_1__0_ cbx_1__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__9_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__9_ccff_tail),
		.chanx_left_out(cbx_1__0__10_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__10_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__10_ccff_tail));

	cbx_1__0_ cbx_1__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__10_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__10_ccff_tail),
		.chanx_left_out(cbx_1__0__11_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__11_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__11_ccff_tail));

	cbx_1__0_ cbx_1__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__11_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__11_ccff_tail),
		.chanx_left_out(cbx_1__0__12_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__12_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__12_ccff_tail));

	cbx_1__0_ cbx_1__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__12_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__12_ccff_tail),
		.chanx_left_out(cbx_1__0__13_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__13_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__13_ccff_tail));

	cbx_1__0_ cbx_1__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__13_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__13_ccff_tail),
		.chanx_left_out(cbx_1__0__14_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__14_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__14_ccff_tail));

	cbx_1__0_ cbx_1__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__14_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__14_ccff_tail),
		.chanx_left_out(cbx_1__0__15_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__15_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__15_ccff_tail));

	cbx_1__0_ cbx_1__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__15_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__15_ccff_tail),
		.chanx_left_out(cbx_1__0__16_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__16_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__16_ccff_tail));

	cbx_1__0_ cbx_1__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__16_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__16_ccff_tail),
		.chanx_left_out(cbx_1__0__17_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__17_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__17_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__18_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__18_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__18_ccff_tail));

	cbx_1__0_ cbx_2__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__17_ccff_tail),
		.chanx_left_out(cbx_1__0__19_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__19_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__19_ccff_tail));

	cbx_1__0_ cbx_2__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__18_ccff_tail),
		.chanx_left_out(cbx_1__0__20_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__20_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__20_ccff_tail));

	cbx_1__0_ cbx_2__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__19_ccff_tail),
		.chanx_left_out(cbx_1__0__21_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__21_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__21_ccff_tail));

	cbx_1__0_ cbx_2__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__20_ccff_tail),
		.chanx_left_out(cbx_1__0__22_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__22_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__22_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__22_ccff_tail));

	cbx_1__0_ cbx_2__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__21_ccff_tail),
		.chanx_left_out(cbx_1__0__23_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__23_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__23_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__23_ccff_tail));

	cbx_1__0_ cbx_2__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__22_ccff_tail),
		.chanx_left_out(cbx_1__0__24_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__24_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__24_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__24_ccff_tail));

	cbx_1__0_ cbx_2__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__23_ccff_tail),
		.chanx_left_out(cbx_1__0__25_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__25_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__25_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__25_ccff_tail));

	cbx_1__0_ cbx_2__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__24_ccff_tail),
		.chanx_left_out(cbx_1__0__26_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__26_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__26_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__26_ccff_tail));

	cbx_1__0_ cbx_2__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__25_ccff_tail),
		.chanx_left_out(cbx_1__0__27_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__27_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__27_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__27_ccff_tail));

	cbx_1__0_ cbx_2__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__26_ccff_tail),
		.chanx_left_out(cbx_1__0__28_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__28_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__28_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__28_ccff_tail));

	cbx_1__0_ cbx_2__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__27_ccff_tail),
		.chanx_left_out(cbx_1__0__29_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__29_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__29_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__29_ccff_tail));

	cbx_1__0_ cbx_2__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__28_ccff_tail),
		.chanx_left_out(cbx_1__0__30_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__30_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__30_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__30_ccff_tail));

	cbx_1__0_ cbx_2__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__29_ccff_tail),
		.chanx_left_out(cbx_1__0__31_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__31_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__31_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__31_ccff_tail));

	cbx_1__0_ cbx_2__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__30_ccff_tail),
		.chanx_left_out(cbx_1__0__32_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__32_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__32_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__32_ccff_tail));

	cbx_1__0_ cbx_2__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__31_ccff_tail),
		.chanx_left_out(cbx_1__0__33_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__33_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__33_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__33_ccff_tail));

	cbx_1__0_ cbx_2__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__32_ccff_tail),
		.chanx_left_out(cbx_1__0__34_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__34_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__34_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__34_ccff_tail));

	cbx_1__0_ cbx_2__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__16_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__33_ccff_tail),
		.chanx_left_out(cbx_1__0__35_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__35_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__35_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__35_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__0__0_chanx_left_out[0:63]),
		.ccff_head(sb_3__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__36_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__36_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__36_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__36_ccff_tail));

	cbx_1__0_ cbx_3__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__17_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__0_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__0_ccff_tail),
		.chanx_left_out(cbx_1__0__37_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__37_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__37_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__37_ccff_tail));

	cbx_1__0_ cbx_3__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__18_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__1_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__1_ccff_tail),
		.chanx_left_out(cbx_1__0__38_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__38_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__38_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__38_ccff_tail));

	cbx_1__0_ cbx_3__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__19_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__2_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__2_ccff_tail),
		.chanx_left_out(cbx_1__0__39_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__39_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__39_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__39_ccff_tail));

	cbx_1__0_ cbx_3__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__20_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__3_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__3_ccff_tail),
		.chanx_left_out(cbx_1__0__40_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__40_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__40_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__40_ccff_tail));

	cbx_1__0_ cbx_3__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__21_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__4_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__4_ccff_tail),
		.chanx_left_out(cbx_1__0__41_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__41_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__41_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__41_ccff_tail));

	cbx_1__0_ cbx_3__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__22_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__5_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__5_ccff_tail),
		.chanx_left_out(cbx_1__0__42_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__42_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__42_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__42_ccff_tail));

	cbx_1__0_ cbx_3__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__23_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__6_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__6_ccff_tail),
		.chanx_left_out(cbx_1__0__43_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__43_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__43_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__43_ccff_tail));

	cbx_1__0_ cbx_3__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__24_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__7_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__7_ccff_tail),
		.chanx_left_out(cbx_1__0__44_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__44_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__44_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__44_ccff_tail));

	cbx_1__0_ cbx_3__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__25_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__8_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__8_ccff_tail),
		.chanx_left_out(cbx_1__0__45_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__45_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__45_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__45_ccff_tail));

	cbx_1__0_ cbx_3__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__26_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__9_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__9_ccff_tail),
		.chanx_left_out(cbx_1__0__46_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__46_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__46_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__46_ccff_tail));

	cbx_1__0_ cbx_3__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__27_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__10_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__10_ccff_tail),
		.chanx_left_out(cbx_1__0__47_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__47_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__47_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__47_ccff_tail));

	cbx_1__0_ cbx_3__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__28_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__11_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__11_ccff_tail),
		.chanx_left_out(cbx_1__0__48_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__48_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__48_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__48_ccff_tail));

	cbx_1__0_ cbx_3__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__29_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__12_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__12_ccff_tail),
		.chanx_left_out(cbx_1__0__49_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__49_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__49_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__49_ccff_tail));

	cbx_1__0_ cbx_3__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__30_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__13_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__13_ccff_tail),
		.chanx_left_out(cbx_1__0__50_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__50_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__50_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__50_ccff_tail));

	cbx_1__0_ cbx_3__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__31_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__14_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__14_ccff_tail),
		.chanx_left_out(cbx_1__0__51_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__51_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__51_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__51_ccff_tail));

	cbx_1__0_ cbx_3__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__32_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__15_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__15_ccff_tail),
		.chanx_left_out(cbx_1__0__52_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__52_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__52_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__52_ccff_tail));

	cbx_1__0_ cbx_3__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__33_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__16_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__16_ccff_tail),
		.chanx_left_out(cbx_1__0__53_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__53_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__53_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__53_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__0__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__54_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__54_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__54_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__54_ccff_tail));

	cbx_1__0_ cbx_5__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__34_ccff_tail),
		.chanx_left_out(cbx_1__0__55_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__55_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__55_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__55_ccff_tail));

	cbx_1__0_ cbx_5__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__35_ccff_tail),
		.chanx_left_out(cbx_1__0__56_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__56_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__56_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__56_ccff_tail));

	cbx_1__0_ cbx_5__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__36_ccff_tail),
		.chanx_left_out(cbx_1__0__57_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__57_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__57_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__57_ccff_tail));

	cbx_1__0_ cbx_5__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__37_ccff_tail),
		.chanx_left_out(cbx_1__0__58_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__58_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__58_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__58_ccff_tail));

	cbx_1__0_ cbx_5__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__38_ccff_tail),
		.chanx_left_out(cbx_1__0__59_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__59_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__59_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__59_ccff_tail));

	cbx_1__0_ cbx_5__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__39_ccff_tail),
		.chanx_left_out(cbx_1__0__60_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__60_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__60_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__60_ccff_tail));

	cbx_1__0_ cbx_5__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__40_ccff_tail),
		.chanx_left_out(cbx_1__0__61_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__61_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__61_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__61_ccff_tail));

	cbx_1__0_ cbx_5__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__41_ccff_tail),
		.chanx_left_out(cbx_1__0__62_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__62_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__62_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__62_ccff_tail));

	cbx_1__0_ cbx_5__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__42_ccff_tail),
		.chanx_left_out(cbx_1__0__63_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__63_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__63_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__63_ccff_tail));

	cbx_1__0_ cbx_5__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__9_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__43_ccff_tail),
		.chanx_left_out(cbx_1__0__64_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__64_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__64_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__64_ccff_tail));

	cbx_1__0_ cbx_5__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__10_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__44_ccff_tail),
		.chanx_left_out(cbx_1__0__65_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__65_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__65_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__65_ccff_tail));

	cbx_1__0_ cbx_5__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__11_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__45_ccff_tail),
		.chanx_left_out(cbx_1__0__66_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__66_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__66_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__66_ccff_tail));

	cbx_1__0_ cbx_5__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__12_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__46_ccff_tail),
		.chanx_left_out(cbx_1__0__67_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__67_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__67_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__67_ccff_tail));

	cbx_1__0_ cbx_5__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__13_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__47_ccff_tail),
		.chanx_left_out(cbx_1__0__68_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__68_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__68_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__68_ccff_tail));

	cbx_1__0_ cbx_5__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__14_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__48_ccff_tail),
		.chanx_left_out(cbx_1__0__69_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__69_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__69_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__69_ccff_tail));

	cbx_1__0_ cbx_5__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__15_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__49_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__49_ccff_tail),
		.chanx_left_out(cbx_1__0__70_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__70_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__70_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__70_ccff_tail));

	cbx_1__0_ cbx_5__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__16_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__50_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__50_ccff_tail),
		.chanx_left_out(cbx_1__0__71_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__71_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__71_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__71_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__72_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__72_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__72_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__72_ccff_tail));

	cbx_1__0_ cbx_6__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__34_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__51_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__51_ccff_tail),
		.chanx_left_out(cbx_1__0__73_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__73_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__73_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__73_ccff_tail));

	cbx_1__0_ cbx_6__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__35_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__52_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__52_ccff_tail),
		.chanx_left_out(cbx_1__0__74_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__74_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__74_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__74_ccff_tail));

	cbx_1__0_ cbx_6__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__36_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__53_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__53_ccff_tail),
		.chanx_left_out(cbx_1__0__75_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__75_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__75_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__75_ccff_tail));

	cbx_1__0_ cbx_6__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__37_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__54_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__54_ccff_tail),
		.chanx_left_out(cbx_1__0__76_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__76_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__76_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__76_ccff_tail));

	cbx_1__0_ cbx_6__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__38_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__55_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__55_ccff_tail),
		.chanx_left_out(cbx_1__0__77_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__77_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__77_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__77_ccff_tail));

	cbx_1__0_ cbx_6__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__39_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__56_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__56_ccff_tail),
		.chanx_left_out(cbx_1__0__78_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__78_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__78_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__78_ccff_tail));

	cbx_1__0_ cbx_6__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__40_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__57_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__57_ccff_tail),
		.chanx_left_out(cbx_1__0__79_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__79_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__79_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__79_ccff_tail));

	cbx_1__0_ cbx_6__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__41_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__58_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__58_ccff_tail),
		.chanx_left_out(cbx_1__0__80_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__80_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__80_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__80_ccff_tail));

	cbx_1__0_ cbx_6__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__42_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__59_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__59_ccff_tail),
		.chanx_left_out(cbx_1__0__81_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__81_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__81_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__81_ccff_tail));

	cbx_1__0_ cbx_6__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__43_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__60_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__60_ccff_tail),
		.chanx_left_out(cbx_1__0__82_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__82_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__82_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__82_ccff_tail));

	cbx_1__0_ cbx_6__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__44_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__61_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__61_ccff_tail),
		.chanx_left_out(cbx_1__0__83_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__83_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__83_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__83_ccff_tail));

	cbx_1__0_ cbx_6__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__45_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__62_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__62_ccff_tail),
		.chanx_left_out(cbx_1__0__84_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__84_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__84_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__84_ccff_tail));

	cbx_1__0_ cbx_6__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__46_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__63_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__63_ccff_tail),
		.chanx_left_out(cbx_1__0__85_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__85_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__85_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__85_ccff_tail));

	cbx_1__0_ cbx_6__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__47_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__64_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__64_ccff_tail),
		.chanx_left_out(cbx_1__0__86_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__86_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__86_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__86_ccff_tail));

	cbx_1__0_ cbx_6__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__48_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__65_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__65_ccff_tail),
		.chanx_left_out(cbx_1__0__87_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__87_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__87_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__87_ccff_tail));

	cbx_1__0_ cbx_6__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__49_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__66_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__66_ccff_tail),
		.chanx_left_out(cbx_1__0__88_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__88_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__88_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__88_ccff_tail));

	cbx_1__0_ cbx_6__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__50_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__67_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__67_ccff_tail),
		.chanx_left_out(cbx_1__0__89_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__89_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__89_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__89_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__90_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__90_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__90_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__90_ccff_tail));

	cbx_1__0_ cbx_7__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__51_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__68_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__68_ccff_tail),
		.chanx_left_out(cbx_1__0__91_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__91_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__91_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__91_ccff_tail));

	cbx_1__0_ cbx_7__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__52_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__69_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__69_ccff_tail),
		.chanx_left_out(cbx_1__0__92_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__92_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__92_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__92_ccff_tail));

	cbx_1__0_ cbx_7__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__53_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__70_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__70_ccff_tail),
		.chanx_left_out(cbx_1__0__93_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__93_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__93_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__93_ccff_tail));

	cbx_1__0_ cbx_7__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__54_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__71_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__71_ccff_tail),
		.chanx_left_out(cbx_1__0__94_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__94_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__94_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__94_ccff_tail));

	cbx_1__0_ cbx_7__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__55_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__72_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__72_ccff_tail),
		.chanx_left_out(cbx_1__0__95_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__95_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__95_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__95_ccff_tail));

	cbx_1__0_ cbx_7__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__56_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__73_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__73_ccff_tail),
		.chanx_left_out(cbx_1__0__96_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__96_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__96_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__96_ccff_tail));

	cbx_1__0_ cbx_7__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__57_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__74_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__74_ccff_tail),
		.chanx_left_out(cbx_1__0__97_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__97_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__97_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__97_ccff_tail));

	cbx_1__0_ cbx_7__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__58_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__75_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__75_ccff_tail),
		.chanx_left_out(cbx_1__0__98_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__98_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__98_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__98_ccff_tail));

	cbx_1__0_ cbx_7__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__59_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__76_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__76_ccff_tail),
		.chanx_left_out(cbx_1__0__99_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__99_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__99_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__99_ccff_tail));

	cbx_1__0_ cbx_7__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__60_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__77_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__77_ccff_tail),
		.chanx_left_out(cbx_1__0__100_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__100_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__100_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__100_ccff_tail));

	cbx_1__0_ cbx_7__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__61_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__78_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__78_ccff_tail),
		.chanx_left_out(cbx_1__0__101_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__101_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__101_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__101_ccff_tail));

	cbx_1__0_ cbx_7__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__62_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__79_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__79_ccff_tail),
		.chanx_left_out(cbx_1__0__102_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__102_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__102_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__102_ccff_tail));

	cbx_1__0_ cbx_7__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__63_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__80_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__80_ccff_tail),
		.chanx_left_out(cbx_1__0__103_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__103_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__103_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__103_ccff_tail));

	cbx_1__0_ cbx_7__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__64_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__81_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__81_ccff_tail),
		.chanx_left_out(cbx_1__0__104_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__104_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__104_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(ccff_tail[9]));

	cbx_1__0_ cbx_7__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__65_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__82_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__82_ccff_tail),
		.chanx_left_out(cbx_1__0__105_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__105_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__105_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__105_ccff_tail));

	cbx_1__0_ cbx_7__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__66_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__83_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__83_ccff_tail),
		.chanx_left_out(cbx_1__0__106_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__106_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__106_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__106_ccff_tail));

	cbx_1__0_ cbx_7__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__67_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__84_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__84_ccff_tail),
		.chanx_left_out(cbx_1__0__107_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__107_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__107_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__107_ccff_tail));

	cbx_1__0_ cbx_8__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__5_ccff_tail),
		.chanx_left_out(cbx_1__0__108_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__108_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__108_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__108_ccff_tail));

	cbx_1__0_ cbx_8__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__68_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__85_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__85_ccff_tail),
		.chanx_left_out(cbx_1__0__109_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__109_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__109_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__109_ccff_tail));

	cbx_1__0_ cbx_8__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__69_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__86_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__86_ccff_tail),
		.chanx_left_out(cbx_1__0__110_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__110_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__110_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__110_ccff_tail));

	cbx_1__0_ cbx_8__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__70_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__87_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__87_ccff_tail),
		.chanx_left_out(cbx_1__0__111_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__111_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__111_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__111_ccff_tail));

	cbx_1__0_ cbx_8__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__71_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__88_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__88_ccff_tail),
		.chanx_left_out(cbx_1__0__112_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__112_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__112_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__112_ccff_tail));

	cbx_1__0_ cbx_8__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__72_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__89_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__89_ccff_tail),
		.chanx_left_out(cbx_1__0__113_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__113_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__113_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__113_ccff_tail));

	cbx_1__0_ cbx_8__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__73_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__90_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__90_ccff_tail),
		.chanx_left_out(cbx_1__0__114_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__114_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__114_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__114_ccff_tail));

	cbx_1__0_ cbx_8__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__74_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__91_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__91_ccff_tail),
		.chanx_left_out(cbx_1__0__115_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__115_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__115_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__115_ccff_tail));

	cbx_1__0_ cbx_8__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__75_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__92_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__92_ccff_tail),
		.chanx_left_out(cbx_1__0__116_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__116_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__116_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__116_ccff_tail));

	cbx_1__0_ cbx_8__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__76_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__93_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__93_ccff_tail),
		.chanx_left_out(cbx_1__0__117_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__117_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__117_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__117_ccff_tail));

	cbx_1__0_ cbx_8__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__77_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__94_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__94_ccff_tail),
		.chanx_left_out(cbx_1__0__118_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__118_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__118_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__118_ccff_tail));

	cbx_1__0_ cbx_8__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__78_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__95_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__95_ccff_tail),
		.chanx_left_out(cbx_1__0__119_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__119_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__119_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__119_ccff_tail));

	cbx_1__0_ cbx_8__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__79_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__96_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__96_ccff_tail),
		.chanx_left_out(cbx_1__0__120_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__120_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__120_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__120_ccff_tail));

	cbx_1__0_ cbx_8__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__80_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__97_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__97_ccff_tail),
		.chanx_left_out(cbx_1__0__121_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__121_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__121_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__121_ccff_tail));

	cbx_1__0_ cbx_8__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__81_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__98_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__98_ccff_tail),
		.chanx_left_out(cbx_1__0__122_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__122_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__122_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__122_ccff_tail));

	cbx_1__0_ cbx_8__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__82_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__99_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__99_ccff_tail),
		.chanx_left_out(cbx_1__0__123_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__123_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__123_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__123_ccff_tail));

	cbx_1__0_ cbx_8__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__83_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__100_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__100_ccff_tail),
		.chanx_left_out(cbx_1__0__124_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__124_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__124_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__124_ccff_tail));

	cbx_1__0_ cbx_8__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__84_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__101_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__101_ccff_tail),
		.chanx_left_out(cbx_1__0__125_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__125_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__125_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__125_ccff_tail));

	cbx_1__0_ cbx_9__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__6_ccff_tail),
		.chanx_left_out(cbx_1__0__126_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__126_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__126_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__126_ccff_tail));

	cbx_1__0_ cbx_9__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__85_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__102_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__102_ccff_tail),
		.chanx_left_out(cbx_1__0__127_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__127_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__127_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__127_ccff_tail));

	cbx_1__0_ cbx_9__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__86_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__103_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__103_ccff_tail),
		.chanx_left_out(cbx_1__0__128_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__128_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__128_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__128_ccff_tail));

	cbx_1__0_ cbx_9__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__87_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__104_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__104_ccff_tail),
		.chanx_left_out(cbx_1__0__129_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__129_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__129_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__129_ccff_tail));

	cbx_1__0_ cbx_9__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__88_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__105_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__105_ccff_tail),
		.chanx_left_out(cbx_1__0__130_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__130_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__130_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__130_ccff_tail));

	cbx_1__0_ cbx_9__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__89_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__106_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__106_ccff_tail),
		.chanx_left_out(cbx_1__0__131_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__131_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__131_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__131_ccff_tail));

	cbx_1__0_ cbx_9__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__90_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__107_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__107_ccff_tail),
		.chanx_left_out(cbx_1__0__132_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__132_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__132_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__132_ccff_tail));

	cbx_1__0_ cbx_9__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__91_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__108_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__108_ccff_tail),
		.chanx_left_out(cbx_1__0__133_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__133_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__133_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__133_ccff_tail));

	cbx_1__0_ cbx_9__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__92_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__109_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__109_ccff_tail),
		.chanx_left_out(cbx_1__0__134_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__134_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__134_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__134_ccff_tail));

	cbx_1__0_ cbx_9__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__93_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__110_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__110_ccff_tail),
		.chanx_left_out(cbx_1__0__135_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__135_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__135_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__135_ccff_tail));

	cbx_1__0_ cbx_9__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__94_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__111_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__111_ccff_tail),
		.chanx_left_out(cbx_1__0__136_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__136_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__136_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__136_ccff_tail));

	cbx_1__0_ cbx_9__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__95_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__112_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__112_ccff_tail),
		.chanx_left_out(cbx_1__0__137_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__137_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__137_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__137_ccff_tail));

	cbx_1__0_ cbx_9__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__96_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__113_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__113_ccff_tail),
		.chanx_left_out(cbx_1__0__138_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__138_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__138_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__138_ccff_tail));

	cbx_1__0_ cbx_9__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__97_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__114_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__114_ccff_tail),
		.chanx_left_out(cbx_1__0__139_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__139_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__139_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__139_ccff_tail));

	cbx_1__0_ cbx_9__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__98_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__115_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__115_ccff_tail),
		.chanx_left_out(cbx_1__0__140_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__140_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__140_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__140_ccff_tail));

	cbx_1__0_ cbx_9__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__99_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__116_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__116_ccff_tail),
		.chanx_left_out(cbx_1__0__141_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__141_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__141_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__141_ccff_tail));

	cbx_1__0_ cbx_9__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__100_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__117_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__117_ccff_tail),
		.chanx_left_out(cbx_1__0__142_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__142_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__142_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__142_ccff_tail));

	cbx_1__0_ cbx_9__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__101_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__118_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__118_ccff_tail),
		.chanx_left_out(cbx_1__0__143_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__143_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__143_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__143_ccff_tail));

	cbx_1__0_ cbx_10__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__0__1_chanx_left_out[0:63]),
		.ccff_head(sb_3__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__144_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__144_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__144_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__144_ccff_tail));

	cbx_1__0_ cbx_10__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__102_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__17_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__17_ccff_tail),
		.chanx_left_out(cbx_1__0__145_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__145_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__145_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__145_ccff_tail));

	cbx_1__0_ cbx_10__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__103_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__18_chanx_left_out[0:63]),
		.ccff_head(ccff_head[3]),
		.chanx_left_out(cbx_1__0__146_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__146_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__146_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__146_ccff_tail));

	cbx_1__0_ cbx_10__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__104_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__19_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__19_ccff_tail),
		.chanx_left_out(cbx_1__0__147_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__147_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__147_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__147_ccff_tail));

	cbx_1__0_ cbx_10__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__105_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__20_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__20_ccff_tail),
		.chanx_left_out(cbx_1__0__148_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__148_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__148_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__148_ccff_tail));

	cbx_1__0_ cbx_10__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__106_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__21_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__21_ccff_tail),
		.chanx_left_out(cbx_1__0__149_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__149_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__149_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__149_ccff_tail));

	cbx_1__0_ cbx_10__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__107_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__22_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__22_ccff_tail),
		.chanx_left_out(cbx_1__0__150_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__150_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__150_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__150_ccff_tail));

	cbx_1__0_ cbx_10__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__108_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__23_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__23_ccff_tail),
		.chanx_left_out(cbx_1__0__151_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__151_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__151_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__151_ccff_tail));

	cbx_1__0_ cbx_10__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__109_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__24_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__24_ccff_tail),
		.chanx_left_out(cbx_1__0__152_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__152_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__152_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__152_ccff_tail));

	cbx_1__0_ cbx_10__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__110_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__25_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__25_ccff_tail),
		.chanx_left_out(cbx_1__0__153_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__153_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__153_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__153_ccff_tail));

	cbx_1__0_ cbx_10__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__111_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__26_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__26_ccff_tail),
		.chanx_left_out(cbx_1__0__154_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__154_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__154_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__154_ccff_tail));

	cbx_1__0_ cbx_10__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__112_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__27_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__27_ccff_tail),
		.chanx_left_out(cbx_1__0__155_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__155_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__155_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__155_ccff_tail));

	cbx_1__0_ cbx_10__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__113_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__28_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__28_ccff_tail),
		.chanx_left_out(cbx_1__0__156_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__156_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__156_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__156_ccff_tail));

	cbx_1__0_ cbx_10__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__114_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__29_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__29_ccff_tail),
		.chanx_left_out(cbx_1__0__157_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__157_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__157_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__157_ccff_tail));

	cbx_1__0_ cbx_10__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__115_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__30_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__30_ccff_tail),
		.chanx_left_out(cbx_1__0__158_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__158_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__158_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__158_ccff_tail));

	cbx_1__0_ cbx_10__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__116_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__31_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__31_ccff_tail),
		.chanx_left_out(cbx_1__0__159_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__159_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__159_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__159_ccff_tail));

	cbx_1__0_ cbx_10__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__117_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__32_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__32_ccff_tail),
		.chanx_left_out(cbx_1__0__160_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__160_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__160_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__160_ccff_tail));

	cbx_1__0_ cbx_10__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__118_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__1__33_chanx_left_out[0:63]),
		.ccff_head(sb_3__1__33_ccff_tail),
		.chanx_left_out(cbx_1__0__161_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__161_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__161_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__161_ccff_tail));

	cbx_1__0_ cbx_12__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__0__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__7_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__7_ccff_tail),
		.chanx_left_out(cbx_1__0__162_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__162_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__162_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__162_ccff_tail));

	cbx_1__0_ cbx_12__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__17_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__119_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__119_ccff_tail),
		.chanx_left_out(cbx_1__0__163_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__163_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__163_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__163_ccff_tail));

	cbx_1__0_ cbx_12__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__18_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__120_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__120_ccff_tail),
		.chanx_left_out(cbx_1__0__164_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__164_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__164_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__164_ccff_tail));

	cbx_1__0_ cbx_12__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__19_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__121_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__121_ccff_tail),
		.chanx_left_out(cbx_1__0__165_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__165_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__165_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__165_ccff_tail));

	cbx_1__0_ cbx_12__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__20_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__122_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__122_ccff_tail),
		.chanx_left_out(cbx_1__0__166_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__166_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__166_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__166_ccff_tail));

	cbx_1__0_ cbx_12__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__21_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__123_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__123_ccff_tail),
		.chanx_left_out(cbx_1__0__167_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__167_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__167_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__167_ccff_tail));

	cbx_1__0_ cbx_12__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__22_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__124_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__124_ccff_tail),
		.chanx_left_out(cbx_1__0__168_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__168_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__168_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__168_ccff_tail));

	cbx_1__0_ cbx_12__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__23_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__125_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__125_ccff_tail),
		.chanx_left_out(cbx_1__0__169_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__169_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__169_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__169_ccff_tail));

	cbx_1__0_ cbx_12__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__24_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__126_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__126_ccff_tail),
		.chanx_left_out(cbx_1__0__170_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__170_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__170_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__170_ccff_tail));

	cbx_1__0_ cbx_12__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__25_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__127_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__127_ccff_tail),
		.chanx_left_out(cbx_1__0__171_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__171_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__171_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__171_ccff_tail));

	cbx_1__0_ cbx_12__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__26_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__128_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__128_ccff_tail),
		.chanx_left_out(cbx_1__0__172_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__172_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__172_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__172_ccff_tail));

	cbx_1__0_ cbx_12__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__27_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__129_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__129_ccff_tail),
		.chanx_left_out(cbx_1__0__173_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__173_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__173_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__173_ccff_tail));

	cbx_1__0_ cbx_12__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__28_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__130_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__130_ccff_tail),
		.chanx_left_out(cbx_1__0__174_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__174_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__174_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__174_ccff_tail));

	cbx_1__0_ cbx_12__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__29_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__131_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__131_ccff_tail),
		.chanx_left_out(cbx_1__0__175_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__175_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__175_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__175_ccff_tail));

	cbx_1__0_ cbx_12__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__30_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__132_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__132_ccff_tail),
		.chanx_left_out(cbx_1__0__176_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__176_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__176_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__176_ccff_tail));

	cbx_1__0_ cbx_12__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__31_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__133_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__133_ccff_tail),
		.chanx_left_out(cbx_1__0__177_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__177_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__177_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__177_ccff_tail));

	cbx_1__0_ cbx_12__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__32_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__134_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__134_ccff_tail),
		.chanx_left_out(cbx_1__0__178_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__178_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__178_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__178_ccff_tail));

	cbx_1__0_ cbx_12__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__1__33_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__135_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__135_ccff_tail),
		.chanx_left_out(cbx_1__0__179_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__179_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__179_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__179_ccff_tail));

	cbx_1__0_ cbx_13__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__0__8_chanx_left_out[0:63]),
		.ccff_head(sb_1__0__8_ccff_tail),
		.chanx_left_out(cbx_1__0__180_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__180_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__180_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__180_ccff_tail));

	cbx_1__0_ cbx_13__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__119_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__136_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__136_ccff_tail),
		.chanx_left_out(cbx_1__0__181_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__181_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__181_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__181_ccff_tail));

	cbx_1__0_ cbx_13__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__120_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__137_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__137_ccff_tail),
		.chanx_left_out(cbx_1__0__182_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__182_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__182_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__182_ccff_tail));

	cbx_1__0_ cbx_13__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__121_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__138_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__138_ccff_tail),
		.chanx_left_out(cbx_1__0__183_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__183_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__183_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__183_ccff_tail));

	cbx_1__0_ cbx_13__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__122_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__139_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__139_ccff_tail),
		.chanx_left_out(cbx_1__0__184_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__184_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__184_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__184_ccff_tail));

	cbx_1__0_ cbx_13__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__123_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__140_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__140_ccff_tail),
		.chanx_left_out(cbx_1__0__185_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__185_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__185_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__185_ccff_tail));

	cbx_1__0_ cbx_13__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__124_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__141_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__141_ccff_tail),
		.chanx_left_out(cbx_1__0__186_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__186_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__186_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__186_ccff_tail));

	cbx_1__0_ cbx_13__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__125_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__142_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__142_ccff_tail),
		.chanx_left_out(cbx_1__0__187_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__187_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__187_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__187_ccff_tail));

	cbx_1__0_ cbx_13__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__126_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__143_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__143_ccff_tail),
		.chanx_left_out(cbx_1__0__188_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__188_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__188_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__188_ccff_tail));

	cbx_1__0_ cbx_13__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__127_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__144_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__144_ccff_tail),
		.chanx_left_out(cbx_1__0__189_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__189_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__189_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__189_ccff_tail));

	cbx_1__0_ cbx_13__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__128_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__145_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__145_ccff_tail),
		.chanx_left_out(cbx_1__0__190_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__190_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__190_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__190_ccff_tail));

	cbx_1__0_ cbx_13__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__129_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__146_chanx_left_out[0:63]),
		.ccff_head(ccff_head[8]),
		.chanx_left_out(cbx_1__0__191_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__191_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__191_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__191_ccff_tail));

	cbx_1__0_ cbx_13__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__130_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__147_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__147_ccff_tail),
		.chanx_left_out(cbx_1__0__192_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__192_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__192_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__192_ccff_tail));

	cbx_1__0_ cbx_13__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__131_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__148_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__148_ccff_tail),
		.chanx_left_out(cbx_1__0__193_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__193_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__193_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__193_ccff_tail));

	cbx_1__0_ cbx_13__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__132_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__149_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__149_ccff_tail),
		.chanx_left_out(cbx_1__0__194_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__194_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__194_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__194_ccff_tail));

	cbx_1__0_ cbx_13__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__133_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__150_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__150_ccff_tail),
		.chanx_left_out(cbx_1__0__195_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__195_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__195_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__195_ccff_tail));

	cbx_1__0_ cbx_13__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__134_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__151_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__151_ccff_tail),
		.chanx_left_out(cbx_1__0__196_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__196_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__196_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__196_ccff_tail));

	cbx_1__0_ cbx_13__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__135_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__1__152_chanx_left_out[0:63]),
		.ccff_head(sb_1__1__152_ccff_tail),
		.chanx_left_out(cbx_1__0__197_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__197_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__197_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__197_ccff_tail));

	cbx_1__0_ cbx_14__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__0__0_chanx_left_out[0:63]),
		.ccff_head(sb_14__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__198_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__198_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__198_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__198_ccff_tail));

	cbx_1__0_ cbx_14__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__136_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__0_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__0_ccff_tail),
		.chanx_left_out(cbx_1__0__199_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__199_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__199_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__199_ccff_tail));

	cbx_1__0_ cbx_14__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__137_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__1_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__1_ccff_tail),
		.chanx_left_out(cbx_1__0__200_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__200_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__200_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__200_ccff_tail));

	cbx_1__0_ cbx_14__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__138_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__2_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__2_ccff_tail),
		.chanx_left_out(cbx_1__0__201_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__201_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__201_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__201_ccff_tail));

	cbx_1__0_ cbx_14__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__139_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__3_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__3_ccff_tail),
		.chanx_left_out(cbx_1__0__202_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__202_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__202_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__202_ccff_tail));

	cbx_1__0_ cbx_14__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__140_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__4_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__4_ccff_tail),
		.chanx_left_out(cbx_1__0__203_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__203_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__203_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__203_ccff_tail));

	cbx_1__0_ cbx_14__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__141_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__5_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__5_ccff_tail),
		.chanx_left_out(cbx_1__0__204_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__204_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__204_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__204_ccff_tail));

	cbx_1__0_ cbx_14__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__142_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__6_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__6_ccff_tail),
		.chanx_left_out(cbx_1__0__205_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__205_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__205_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__205_ccff_tail));

	cbx_1__0_ cbx_14__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__143_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__7_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__7_ccff_tail),
		.chanx_left_out(cbx_1__0__206_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__206_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__206_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__206_ccff_tail));

	cbx_1__0_ cbx_14__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__144_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__8_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__8_ccff_tail),
		.chanx_left_out(cbx_1__0__207_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__207_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__207_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__207_ccff_tail));

	cbx_1__0_ cbx_14__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__145_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__9_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__9_ccff_tail),
		.chanx_left_out(cbx_1__0__208_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__208_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__208_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__208_ccff_tail));

	cbx_1__0_ cbx_14__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__146_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__10_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__10_ccff_tail),
		.chanx_left_out(cbx_1__0__209_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__209_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__209_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__209_ccff_tail));

	cbx_1__0_ cbx_14__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__147_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__11_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__11_ccff_tail),
		.chanx_left_out(cbx_1__0__210_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__210_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__210_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__210_ccff_tail));

	cbx_1__0_ cbx_14__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__148_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__12_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__12_ccff_tail),
		.chanx_left_out(cbx_1__0__211_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__211_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__211_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__211_ccff_tail));

	cbx_1__0_ cbx_14__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__149_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__13_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__13_ccff_tail),
		.chanx_left_out(cbx_1__0__212_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__212_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__212_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__212_ccff_tail));

	cbx_1__0_ cbx_14__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__150_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__14_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__14_ccff_tail),
		.chanx_left_out(cbx_1__0__213_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__213_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__213_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__213_ccff_tail));

	cbx_1__0_ cbx_14__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__151_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__15_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__15_ccff_tail),
		.chanx_left_out(cbx_1__0__214_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__214_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__214_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__214_ccff_tail));

	cbx_1__0_ cbx_14__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__152_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__1__16_chanx_left_out[0:63]),
		.ccff_head(sb_14__1__16_ccff_tail),
		.chanx_left_out(cbx_1__0__215_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__0__215_chanx_right_out[0:63]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__215_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__215_ccff_tail));

	cbx_1__18_ cbx_1__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__18__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__0_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__0_ccff_tail),
		.chanx_left_out(cbx_1__18__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__0_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__0_ccff_tail));

	cbx_1__18_ cbx_2__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__1_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__1_ccff_tail),
		.chanx_left_out(cbx_1__18__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__1_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__1_ccff_tail));

	cbx_1__18_ cbx_3__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__18__0_chanx_left_out[0:63]),
		.ccff_head(sb_3__18__0_ccff_tail),
		.chanx_left_out(cbx_1__18__2_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__2_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__2_ccff_tail));

	cbx_1__18_ cbx_5__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__18__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__2_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__2_ccff_tail),
		.chanx_left_out(cbx_1__18__3_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__3_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__3_ccff_tail));

	cbx_1__18_ cbx_6__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__3_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__3_ccff_tail),
		.chanx_left_out(cbx_1__18__4_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__4_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__4_ccff_tail));

	cbx_1__18_ cbx_7__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__4_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__4_ccff_tail),
		.chanx_left_out(cbx_1__18__5_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__5_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__5_ccff_tail));

	cbx_1__18_ cbx_8__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__5_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__5_ccff_tail),
		.chanx_left_out(cbx_1__18__6_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__6_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__6_ccff_tail));

	cbx_1__18_ cbx_9__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__6_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__6_ccff_tail),
		.chanx_left_out(cbx_1__18__7_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__7_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__7_ccff_tail));

	cbx_1__18_ cbx_10__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_3__18__1_chanx_left_out[0:63]),
		.ccff_head(sb_3__18__1_ccff_tail),
		.chanx_left_out(cbx_1__18__8_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__8_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__8_ccff_tail));

	cbx_1__18_ cbx_12__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__18__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__7_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__7_ccff_tail),
		.chanx_left_out(cbx_1__18__9_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__9_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__9_ccff_tail));

	cbx_1__18_ cbx_13__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_1__18__8_chanx_left_out[0:63]),
		.ccff_head(sb_1__18__8_ccff_tail),
		.chanx_left_out(cbx_1__18__10_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__10_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__10_ccff_tail));

	cbx_1__18_ cbx_14__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__18__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_14__18__0_chanx_left_out[0:63]),
		.ccff_head(sb_14__18__0_ccff_tail),
		.chanx_left_out(cbx_1__18__11_chanx_left_out[0:63]),
		.chanx_right_out(cbx_1__18__11_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__18__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__18__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__18__11_ccff_tail));

	cbx_4__0_ cbx_4__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__0__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__0__0_chanx_left_out[0:63]),
		.ccff_head(sb_4__0__0_ccff_tail),
		.chanx_left_out(cbx_4__0__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__0__0_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_4__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_4__0__0_ccff_tail));

	cbx_4__0_ cbx_11__0_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__0__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__0__1_chanx_left_out[0:63]),
		.ccff_head(sb_4__0__1_ccff_tail),
		.chanx_left_out(cbx_4__0__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__0__1_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_4__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_4__0__1_ccff_tail));

	cbx_4__1_ cbx_4__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__0_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__0_ccff_tail),
		.chanx_left_out(cbx_4__1__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__0_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__0_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__0_ccff_tail));

	cbx_4__1_ cbx_4__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__2_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__2_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__2_ccff_tail),
		.chanx_left_out(cbx_4__1__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__1_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__1_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__1_ccff_tail));

	cbx_4__1_ cbx_4__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__4_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__4_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__4_ccff_tail),
		.chanx_left_out(cbx_4__1__2_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__2_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__2_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__2_ccff_tail));

	cbx_4__1_ cbx_4__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__6_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__6_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__6_ccff_tail),
		.chanx_left_out(cbx_4__1__3_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__3_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__3_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__3_ccff_tail));

	cbx_4__1_ cbx_4__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__8_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__8_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__8_ccff_tail),
		.chanx_left_out(cbx_4__1__4_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__4_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__4_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__4_ccff_tail));

	cbx_4__1_ cbx_4__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__10_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__10_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__10_ccff_tail),
		.chanx_left_out(cbx_4__1__5_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__5_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__5_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__5_ccff_tail));

	cbx_4__1_ cbx_4__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__12_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__12_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__12_ccff_tail),
		.chanx_left_out(cbx_4__1__6_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__6_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__6_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__6_ccff_tail));

	cbx_4__1_ cbx_4__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__14_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__14_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__14_ccff_tail),
		.chanx_left_out(cbx_4__1__7_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__7_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__7_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__7_ccff_tail));

	cbx_4__1_ cbx_4__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__16_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__16_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__16_ccff_tail),
		.chanx_left_out(cbx_4__1__8_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__8_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__8_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__8_ccff_tail));

	cbx_4__1_ cbx_11__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__17_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__17_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__17_ccff_tail),
		.chanx_left_out(cbx_4__1__9_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__9_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__9_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__9_ccff_tail));

	cbx_4__1_ cbx_11__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__19_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__19_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__19_ccff_tail),
		.chanx_left_out(cbx_4__1__10_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__10_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__10_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__10_ccff_tail));

	cbx_4__1_ cbx_11__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__21_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__21_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__21_ccff_tail),
		.chanx_left_out(cbx_4__1__11_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__11_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__11_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__11_ccff_tail));

	cbx_4__1_ cbx_11__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__23_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__23_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__23_ccff_tail),
		.chanx_left_out(cbx_4__1__12_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__12_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__12_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__12_ccff_tail));

	cbx_4__1_ cbx_11__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__25_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__25_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__25_ccff_tail),
		.chanx_left_out(cbx_4__1__13_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__13_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__13_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__13_ccff_tail));

	cbx_4__1_ cbx_11__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__27_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__27_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__27_ccff_tail),
		.chanx_left_out(cbx_4__1__14_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__14_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__14_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__14_ccff_tail));

	cbx_4__1_ cbx_11__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__29_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__29_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__29_ccff_tail),
		.chanx_left_out(cbx_4__1__15_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__15_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__15_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__15_ccff_tail));

	cbx_4__1_ cbx_11__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__31_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__31_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__31_ccff_tail),
		.chanx_left_out(cbx_4__1__16_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__16_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__16_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__16_ccff_tail));

	cbx_4__1_ cbx_11__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__33_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__33_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__33_ccff_tail),
		.chanx_left_out(cbx_4__1__17_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__1__17_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_raddr_4_),
		.top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_(cbx_4__1__17_top_grid_bottom_width_0_height_1_subtile_0__pin_data_in_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_(cbx_4__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_data_in_6_),
		.ccff_tail(cbx_4__1__17_ccff_tail));

	cbx_4__2_ cbx_4__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__1_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__1_ccff_tail),
		.chanx_left_out(cbx_4__2__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__0_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__0_ccff_tail));

	cbx_4__2_ cbx_4__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__3_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__3_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__3_ccff_tail),
		.chanx_left_out(cbx_4__2__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__1_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__1_ccff_tail));

	cbx_4__2_ cbx_4__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__5_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__5_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__5_ccff_tail),
		.chanx_left_out(cbx_4__2__2_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__2_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__2_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__2_ccff_tail));

	cbx_4__2_ cbx_4__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__7_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__7_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__7_ccff_tail),
		.chanx_left_out(cbx_4__2__3_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__3_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__3_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__3_ccff_tail));

	cbx_4__2_ cbx_4__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__9_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__9_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__9_ccff_tail),
		.chanx_left_out(cbx_4__2__4_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__4_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__4_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__4_ccff_tail));

	cbx_4__2_ cbx_4__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__11_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__11_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__11_ccff_tail),
		.chanx_left_out(cbx_4__2__5_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__5_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__5_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__5_ccff_tail));

	cbx_4__2_ cbx_4__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__13_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__13_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__13_ccff_tail),
		.chanx_left_out(cbx_4__2__6_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__6_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__6_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__6_ccff_tail));

	cbx_4__2_ cbx_4__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__15_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__15_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__15_ccff_tail),
		.chanx_left_out(cbx_4__2__7_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__7_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__7_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__7_ccff_tail));

	cbx_4__2_ cbx_11__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__18_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__18_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__18_ccff_tail),
		.chanx_left_out(cbx_4__2__8_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__8_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__8_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__8_ccff_tail));

	cbx_4__2_ cbx_11__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__20_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__20_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__20_ccff_tail),
		.chanx_left_out(cbx_4__2__9_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__9_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__9_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__9_ccff_tail));

	cbx_4__2_ cbx_11__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__22_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__22_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__22_ccff_tail),
		.chanx_left_out(cbx_4__2__10_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__10_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__10_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__10_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__10_ccff_tail));

	cbx_4__2_ cbx_11__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__24_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__24_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__24_ccff_tail),
		.chanx_left_out(cbx_4__2__11_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__11_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__11_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__11_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__11_ccff_tail));

	cbx_4__2_ cbx_11__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__26_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__26_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__26_ccff_tail),
		.chanx_left_out(cbx_4__2__12_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__12_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__12_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__12_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__12_ccff_tail));

	cbx_4__2_ cbx_11__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__28_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__28_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__28_ccff_tail),
		.chanx_left_out(cbx_4__2__13_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__13_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__13_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__13_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__13_ccff_tail));

	cbx_4__2_ cbx_11__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__30_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__30_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__30_ccff_tail),
		.chanx_left_out(cbx_4__2__14_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__14_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__14_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__14_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__14_ccff_tail));

	cbx_4__2_ cbx_11__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__32_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__1__32_chanx_left_out[0:63]),
		.ccff_head(sb_4__1__32_ccff_tail),
		.chanx_left_out(cbx_4__2__15_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__2__15_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_(cbx_4__2__15_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_2_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__2__15_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__2__15_ccff_tail));

	cbx_4__18_ cbx_4__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__18__0_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__18__0_chanx_left_out[0:63]),
		.ccff_head(sb_4__18__0_ccff_tail),
		.chanx_left_out(cbx_4__18__0_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__18__0_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__18__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__18__0_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__18__0_ccff_tail));

	cbx_4__18_ cbx_11__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__18__1_chanx_right_out[0:63]),
		.chanx_right_in(sb_4__18__1_chanx_left_out[0:63]),
		.ccff_head(sb_4__18__1_ccff_tail),
		.chanx_left_out(cbx_4__18__1_chanx_left_out[0:63]),
		.chanx_right_out(cbx_4__18__1_chanx_right_out[0:63]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__18__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_waddr_1_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_0_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_raddr_8_),
		.bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_(cbx_4__18__1_bottom_grid_top_width_0_height_1_subtile_0__pin_data_in_7_),
		.ccff_tail(cbx_4__18__1_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:63]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__4_ccff_tail),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__5_ccff_tail));

	cby_0__1_ cby_0__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__5_ccff_tail),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__6_ccff_tail));

	cby_0__1_ cby_0__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__7_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__6_ccff_tail),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__7_ccff_tail));

	cby_0__1_ cby_0__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__7_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__8_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__7_ccff_tail),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__8_ccff_tail));

	cby_0__1_ cby_0__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__8_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__9_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__8_ccff_tail),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__9_ccff_tail));

	cby_0__1_ cby_0__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__9_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__10_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__9_ccff_tail),
		.chany_bottom_out(cby_0__1__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__10_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__10_ccff_tail));

	cby_0__1_ cby_0__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__10_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__11_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__10_ccff_tail),
		.chany_bottom_out(cby_0__1__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__11_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__11_ccff_tail));

	cby_0__1_ cby_0__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__11_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__12_chany_bottom_out[0:63]),
		.ccff_head(ccff_head[1]),
		.chany_bottom_out(cby_0__1__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__12_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__12_ccff_tail));

	cby_0__1_ cby_0__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__12_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__13_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__12_ccff_tail),
		.chany_bottom_out(cby_0__1__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__13_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__13_ccff_tail));

	cby_0__1_ cby_0__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__13_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__14_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__13_ccff_tail),
		.chany_bottom_out(cby_0__1__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__14_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__14_ccff_tail));

	cby_0__1_ cby_0__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__14_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__15_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__14_ccff_tail),
		.chany_bottom_out(cby_0__1__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__15_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__15_ccff_tail));

	cby_0__1_ cby_0__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__15_chany_top_out[0:63]),
		.chany_top_in(sb_0__1__16_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__15_ccff_tail),
		.chany_bottom_out(cby_0__1__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__16_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__16_ccff_tail));

	cby_0__1_ cby_0__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__16_chany_top_out[0:63]),
		.chany_top_in(sb_0__18__0_chany_bottom_out[0:63]),
		.ccff_head(sb_0__1__16_ccff_tail),
		.chany_bottom_out(cby_0__1__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_0__1__17_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__17_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_1__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_1__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_1__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:63]),
		.ccff_head(ccff_head[5]),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_1__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__7_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_1__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__8_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_1__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__9_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_1__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__10_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_1__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__11_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_1__1_ cby_1__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__12_ccff_tail),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__12_ccff_tail));

	cby_1__1_ cby_1__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__13_ccff_tail),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__13_ccff_tail));

	cby_1__1_ cby_1__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__14_ccff_tail),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__14_ccff_tail));

	cby_1__1_ cby_1__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__15_ccff_tail),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__15_ccff_tail));

	cby_1__1_ cby_1__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__16_ccff_tail),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__16_ccff_tail));

	cby_1__1_ cby_1__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__16_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__17_ccff_tail),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__17_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__18_ccff_tail),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__18_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__17_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__19_ccff_tail),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__19_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__18_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__20_ccff_tail),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__20_ccff_tail));

	cby_1__1_ cby_2__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__19_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__21_ccff_tail),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__21_ccff_tail));

	cby_1__1_ cby_2__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__20_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__22_ccff_tail),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__22_ccff_tail));

	cby_1__1_ cby_2__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__21_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__23_ccff_tail),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__23_ccff_tail));

	cby_1__1_ cby_2__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__22_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__24_ccff_tail),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__24_ccff_tail));

	cby_1__1_ cby_2__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__23_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__25_ccff_tail),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__25_ccff_tail));

	cby_1__1_ cby_2__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__24_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__26_ccff_tail),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__26_ccff_tail));

	cby_1__1_ cby_2__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__25_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__27_ccff_tail),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__27_ccff_tail));

	cby_1__1_ cby_2__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__26_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__28_ccff_tail),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__28_ccff_tail));

	cby_1__1_ cby_2__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__27_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__29_ccff_tail),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__29_ccff_tail));

	cby_1__1_ cby_2__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__28_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__30_ccff_tail),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__30_ccff_tail));

	cby_1__1_ cby_2__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__29_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__31_ccff_tail),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__31_ccff_tail));

	cby_1__1_ cby_2__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__30_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__32_ccff_tail),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__32_ccff_tail));

	cby_1__1_ cby_2__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__31_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__33_ccff_tail),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__33_ccff_tail));

	cby_1__1_ cby_2__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__32_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__34_ccff_tail),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__34_ccff_tail));

	cby_1__1_ cby_2__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__33_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__35_ccff_tail),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__35_ccff_tail));

	cby_1__1_ cby_5__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__54_ccff_tail),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__36_ccff_tail));

	cby_1__1_ cby_5__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__34_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__55_ccff_tail),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__37_ccff_tail));

	cby_1__1_ cby_5__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__35_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__56_ccff_tail),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__38_ccff_tail));

	cby_1__1_ cby_5__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__36_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__57_ccff_tail),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__39_ccff_tail));

	cby_1__1_ cby_5__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__37_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__58_ccff_tail),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__40_ccff_tail));

	cby_1__1_ cby_5__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__38_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__59_ccff_tail),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__41_ccff_tail));

	cby_1__1_ cby_5__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__39_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__60_ccff_tail),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__42_ccff_tail));

	cby_1__1_ cby_5__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__40_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__61_ccff_tail),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__43_ccff_tail));

	cby_1__1_ cby_5__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__41_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__62_ccff_tail),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__44_ccff_tail));

	cby_1__1_ cby_5__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__42_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__63_ccff_tail),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__45_ccff_tail));

	cby_1__1_ cby_5__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__43_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__64_ccff_tail),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__46_ccff_tail));

	cby_1__1_ cby_5__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__44_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__65_ccff_tail),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__47_ccff_tail));

	cby_1__1_ cby_5__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__45_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__66_ccff_tail),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__48_ccff_tail));

	cby_1__1_ cby_5__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__46_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__67_ccff_tail),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__49_ccff_tail));

	cby_1__1_ cby_5__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__47_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__68_ccff_tail),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__50_ccff_tail));

	cby_1__1_ cby_5__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__48_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__49_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__69_ccff_tail),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__51_ccff_tail));

	cby_1__1_ cby_5__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__49_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__50_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__70_ccff_tail),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__52_ccff_tail));

	cby_1__1_ cby_5__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__50_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__2_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__71_ccff_tail),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__53_ccff_tail));

	cby_1__1_ cby_6__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__51_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__72_ccff_tail),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__54_ccff_tail));

	cby_1__1_ cby_6__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__51_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__52_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__73_ccff_tail),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__55_ccff_tail));

	cby_1__1_ cby_6__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__52_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__53_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__74_ccff_tail),
		.chany_bottom_out(cby_1__1__56_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__56_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__56_ccff_tail));

	cby_1__1_ cby_6__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__53_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__54_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__75_ccff_tail),
		.chany_bottom_out(cby_1__1__57_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__57_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__57_ccff_tail));

	cby_1__1_ cby_6__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__54_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__55_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__76_ccff_tail),
		.chany_bottom_out(cby_1__1__58_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__58_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__58_ccff_tail));

	cby_1__1_ cby_6__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__55_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__56_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__77_ccff_tail),
		.chany_bottom_out(cby_1__1__59_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__59_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__59_ccff_tail));

	cby_1__1_ cby_6__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__56_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__57_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__78_ccff_tail),
		.chany_bottom_out(cby_1__1__60_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__60_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__60_ccff_tail));

	cby_1__1_ cby_6__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__57_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__58_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__79_ccff_tail),
		.chany_bottom_out(cby_1__1__61_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__61_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__61_ccff_tail));

	cby_1__1_ cby_6__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__58_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__59_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__80_ccff_tail),
		.chany_bottom_out(cby_1__1__62_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__62_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__62_ccff_tail));

	cby_1__1_ cby_6__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__59_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__60_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__81_ccff_tail),
		.chany_bottom_out(cby_1__1__63_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__63_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__63_ccff_tail));

	cby_1__1_ cby_6__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__60_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__61_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__82_ccff_tail),
		.chany_bottom_out(cby_1__1__64_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__64_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__64_ccff_tail));

	cby_1__1_ cby_6__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__61_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__62_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__83_ccff_tail),
		.chany_bottom_out(cby_1__1__65_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__65_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__65_ccff_tail));

	cby_1__1_ cby_6__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__62_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__63_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__84_ccff_tail),
		.chany_bottom_out(cby_1__1__66_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__66_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__66_ccff_tail));

	cby_1__1_ cby_6__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__63_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__64_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__85_ccff_tail),
		.chany_bottom_out(cby_1__1__67_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__67_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__67_ccff_tail));

	cby_1__1_ cby_6__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__64_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__65_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__86_ccff_tail),
		.chany_bottom_out(cby_1__1__68_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__68_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__68_ccff_tail));

	cby_1__1_ cby_6__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__65_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__66_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__87_ccff_tail),
		.chany_bottom_out(cby_1__1__69_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__69_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__69_ccff_tail));

	cby_1__1_ cby_6__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__66_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__67_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__88_ccff_tail),
		.chany_bottom_out(cby_1__1__70_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__70_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__70_ccff_tail));

	cby_1__1_ cby_6__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__67_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__3_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__89_ccff_tail),
		.chany_bottom_out(cby_1__1__71_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__71_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__71_ccff_tail));

	cby_1__1_ cby_7__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__68_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__90_ccff_tail),
		.chany_bottom_out(cby_1__1__72_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__72_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__72_ccff_tail));

	cby_1__1_ cby_7__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__68_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__69_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__91_ccff_tail),
		.chany_bottom_out(cby_1__1__73_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__73_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__73_ccff_tail));

	cby_1__1_ cby_7__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__69_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__70_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__92_ccff_tail),
		.chany_bottom_out(cby_1__1__74_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__74_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__74_ccff_tail));

	cby_1__1_ cby_7__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__70_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__71_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__93_ccff_tail),
		.chany_bottom_out(cby_1__1__75_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__75_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__75_ccff_tail));

	cby_1__1_ cby_7__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__71_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__72_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__94_ccff_tail),
		.chany_bottom_out(cby_1__1__76_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__76_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__76_ccff_tail));

	cby_1__1_ cby_7__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__72_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__73_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__95_ccff_tail),
		.chany_bottom_out(cby_1__1__77_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__77_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__77_ccff_tail));

	cby_1__1_ cby_7__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__73_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__74_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__96_ccff_tail),
		.chany_bottom_out(cby_1__1__78_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__78_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__78_ccff_tail));

	cby_1__1_ cby_7__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__74_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__75_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__97_ccff_tail),
		.chany_bottom_out(cby_1__1__79_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__79_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__79_ccff_tail));

	cby_1__1_ cby_7__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__75_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__76_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__98_ccff_tail),
		.chany_bottom_out(cby_1__1__80_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__80_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__80_ccff_tail));

	cby_1__1_ cby_7__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__76_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__77_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__99_ccff_tail),
		.chany_bottom_out(cby_1__1__81_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__81_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__81_ccff_tail));

	cby_1__1_ cby_7__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__77_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__78_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__100_ccff_tail),
		.chany_bottom_out(cby_1__1__82_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__82_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__82_ccff_tail));

	cby_1__1_ cby_7__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__78_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__79_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__101_ccff_tail),
		.chany_bottom_out(cby_1__1__83_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__83_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__83_ccff_tail));

	cby_1__1_ cby_7__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__79_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__80_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__102_ccff_tail),
		.chany_bottom_out(cby_1__1__84_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__84_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__84_ccff_tail));

	cby_1__1_ cby_7__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__80_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__81_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__103_ccff_tail),
		.chany_bottom_out(cby_1__1__85_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__85_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__85_ccff_tail));

	cby_1__1_ cby_7__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__81_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__82_chany_bottom_out[0:63]),
		.ccff_head(ccff_head[10]),
		.chany_bottom_out(cby_1__1__86_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__86_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__86_ccff_tail));

	cby_1__1_ cby_7__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__82_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__83_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__105_ccff_tail),
		.chany_bottom_out(cby_1__1__87_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__87_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__87_ccff_tail));

	cby_1__1_ cby_7__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__83_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__84_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__106_ccff_tail),
		.chany_bottom_out(cby_1__1__88_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__88_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__88_ccff_tail));

	cby_1__1_ cby_7__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__84_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__4_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__107_ccff_tail),
		.chany_bottom_out(cby_1__1__89_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__89_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__89_ccff_tail));

	cby_1__1_ cby_8__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__85_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__108_ccff_tail),
		.chany_bottom_out(cby_1__1__90_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__90_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__90_ccff_tail));

	cby_1__1_ cby_8__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__85_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__86_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__109_ccff_tail),
		.chany_bottom_out(cby_1__1__91_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__91_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__91_ccff_tail));

	cby_1__1_ cby_8__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__86_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__87_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__110_ccff_tail),
		.chany_bottom_out(cby_1__1__92_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__92_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__92_ccff_tail));

	cby_1__1_ cby_8__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__87_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__88_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__111_ccff_tail),
		.chany_bottom_out(cby_1__1__93_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__93_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__93_ccff_tail));

	cby_1__1_ cby_8__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__88_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__89_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__112_ccff_tail),
		.chany_bottom_out(cby_1__1__94_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__94_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__94_ccff_tail));

	cby_1__1_ cby_8__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__89_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__90_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__113_ccff_tail),
		.chany_bottom_out(cby_1__1__95_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__95_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__95_ccff_tail));

	cby_1__1_ cby_8__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__90_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__91_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__114_ccff_tail),
		.chany_bottom_out(cby_1__1__96_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__96_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__96_ccff_tail));

	cby_1__1_ cby_8__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__91_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__92_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__115_ccff_tail),
		.chany_bottom_out(cby_1__1__97_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__97_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__97_ccff_tail));

	cby_1__1_ cby_8__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__92_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__93_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__116_ccff_tail),
		.chany_bottom_out(cby_1__1__98_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__98_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__98_ccff_tail));

	cby_1__1_ cby_8__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__93_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__94_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__117_ccff_tail),
		.chany_bottom_out(cby_1__1__99_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__99_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__99_ccff_tail));

	cby_1__1_ cby_8__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__94_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__95_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__118_ccff_tail),
		.chany_bottom_out(cby_1__1__100_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__100_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__100_ccff_tail));

	cby_1__1_ cby_8__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__95_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__96_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__119_ccff_tail),
		.chany_bottom_out(cby_1__1__101_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__101_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__101_ccff_tail));

	cby_1__1_ cby_8__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__96_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__97_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__120_ccff_tail),
		.chany_bottom_out(cby_1__1__102_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__102_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__102_ccff_tail));

	cby_1__1_ cby_8__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__97_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__98_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__121_ccff_tail),
		.chany_bottom_out(cby_1__1__103_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__103_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__103_ccff_tail));

	cby_1__1_ cby_8__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__98_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__99_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__122_ccff_tail),
		.chany_bottom_out(cby_1__1__104_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__104_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__104_ccff_tail));

	cby_1__1_ cby_8__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__99_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__100_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__123_ccff_tail),
		.chany_bottom_out(cby_1__1__105_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__105_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__105_ccff_tail));

	cby_1__1_ cby_8__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__100_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__101_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__124_ccff_tail),
		.chany_bottom_out(cby_1__1__106_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__106_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__106_ccff_tail));

	cby_1__1_ cby_8__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__101_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__5_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__125_ccff_tail),
		.chany_bottom_out(cby_1__1__107_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__107_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__107_ccff_tail));

	cby_1__1_ cby_9__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__102_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__126_ccff_tail),
		.chany_bottom_out(cby_1__1__108_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__108_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__108_ccff_tail));

	cby_1__1_ cby_9__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__102_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__103_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__127_ccff_tail),
		.chany_bottom_out(cby_1__1__109_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__109_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__109_ccff_tail));

	cby_1__1_ cby_9__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__103_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__104_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__128_ccff_tail),
		.chany_bottom_out(cby_1__1__110_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__110_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__110_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__110_ccff_tail));

	cby_1__1_ cby_9__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__104_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__105_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__129_ccff_tail),
		.chany_bottom_out(cby_1__1__111_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__111_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__111_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__111_ccff_tail));

	cby_1__1_ cby_9__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__105_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__106_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__130_ccff_tail),
		.chany_bottom_out(cby_1__1__112_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__112_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__112_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__112_ccff_tail));

	cby_1__1_ cby_9__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__106_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__107_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__131_ccff_tail),
		.chany_bottom_out(cby_1__1__113_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__113_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__113_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__113_ccff_tail));

	cby_1__1_ cby_9__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__107_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__108_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__132_ccff_tail),
		.chany_bottom_out(cby_1__1__114_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__114_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__114_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__114_ccff_tail));

	cby_1__1_ cby_9__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__108_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__109_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__133_ccff_tail),
		.chany_bottom_out(cby_1__1__115_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__115_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__115_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__115_ccff_tail));

	cby_1__1_ cby_9__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__109_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__110_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__134_ccff_tail),
		.chany_bottom_out(cby_1__1__116_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__116_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__116_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__116_ccff_tail));

	cby_1__1_ cby_9__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__110_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__111_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__135_ccff_tail),
		.chany_bottom_out(cby_1__1__117_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__117_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__117_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(ccff_tail[6]));

	cby_1__1_ cby_9__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__111_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__112_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__136_ccff_tail),
		.chany_bottom_out(cby_1__1__118_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__118_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__118_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__118_ccff_tail));

	cby_1__1_ cby_9__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__112_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__113_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__137_ccff_tail),
		.chany_bottom_out(cby_1__1__119_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__119_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__119_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__119_ccff_tail));

	cby_1__1_ cby_9__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__113_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__114_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__138_ccff_tail),
		.chany_bottom_out(cby_1__1__120_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__120_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__120_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__120_ccff_tail));

	cby_1__1_ cby_9__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__114_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__115_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__139_ccff_tail),
		.chany_bottom_out(cby_1__1__121_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__121_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__121_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__121_ccff_tail));

	cby_1__1_ cby_9__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__115_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__116_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__140_ccff_tail),
		.chany_bottom_out(cby_1__1__122_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__122_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__122_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__122_ccff_tail));

	cby_1__1_ cby_9__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__116_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__117_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__141_ccff_tail),
		.chany_bottom_out(cby_1__1__123_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__123_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__123_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__123_ccff_tail));

	cby_1__1_ cby_9__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__117_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__118_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__142_ccff_tail),
		.chany_bottom_out(cby_1__1__124_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__124_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__124_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__124_ccff_tail));

	cby_1__1_ cby_9__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__118_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__6_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__143_ccff_tail),
		.chany_bottom_out(cby_1__1__125_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__125_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__125_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__125_ccff_tail));

	cby_1__1_ cby_12__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__7_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__119_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__162_ccff_tail),
		.chany_bottom_out(cby_1__1__126_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__126_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__126_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__126_ccff_tail));

	cby_1__1_ cby_12__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__119_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__120_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__163_ccff_tail),
		.chany_bottom_out(cby_1__1__127_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__127_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__127_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__127_ccff_tail));

	cby_1__1_ cby_12__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__120_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__121_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__164_ccff_tail),
		.chany_bottom_out(cby_1__1__128_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__128_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__128_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__128_ccff_tail));

	cby_1__1_ cby_12__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__121_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__122_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__165_ccff_tail),
		.chany_bottom_out(cby_1__1__129_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__129_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__129_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__129_ccff_tail));

	cby_1__1_ cby_12__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__122_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__123_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__166_ccff_tail),
		.chany_bottom_out(cby_1__1__130_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__130_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__130_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__130_ccff_tail));

	cby_1__1_ cby_12__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__123_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__124_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__167_ccff_tail),
		.chany_bottom_out(cby_1__1__131_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__131_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__131_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__131_ccff_tail));

	cby_1__1_ cby_12__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__124_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__125_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__168_ccff_tail),
		.chany_bottom_out(cby_1__1__132_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__132_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__132_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__132_ccff_tail));

	cby_1__1_ cby_12__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__125_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__126_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__169_ccff_tail),
		.chany_bottom_out(cby_1__1__133_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__133_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__133_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__133_ccff_tail));

	cby_1__1_ cby_12__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__126_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__127_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__170_ccff_tail),
		.chany_bottom_out(cby_1__1__134_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__134_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__134_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__134_ccff_tail));

	cby_1__1_ cby_12__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__127_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__128_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__171_ccff_tail),
		.chany_bottom_out(cby_1__1__135_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__135_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__135_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__135_ccff_tail));

	cby_1__1_ cby_12__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__128_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__129_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__172_ccff_tail),
		.chany_bottom_out(cby_1__1__136_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__136_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__136_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__136_ccff_tail));

	cby_1__1_ cby_12__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__129_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__130_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__173_ccff_tail),
		.chany_bottom_out(cby_1__1__137_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__137_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__137_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__137_ccff_tail));

	cby_1__1_ cby_12__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__130_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__131_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__174_ccff_tail),
		.chany_bottom_out(cby_1__1__138_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__138_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__138_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__138_ccff_tail));

	cby_1__1_ cby_12__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__131_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__132_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__175_ccff_tail),
		.chany_bottom_out(cby_1__1__139_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__139_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__139_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__139_ccff_tail));

	cby_1__1_ cby_12__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__132_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__133_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__176_ccff_tail),
		.chany_bottom_out(cby_1__1__140_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__140_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__140_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__140_ccff_tail));

	cby_1__1_ cby_12__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__133_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__134_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__177_ccff_tail),
		.chany_bottom_out(cby_1__1__141_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__141_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__141_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__141_ccff_tail));

	cby_1__1_ cby_12__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__134_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__135_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__178_ccff_tail),
		.chany_bottom_out(cby_1__1__142_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__142_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__142_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__142_ccff_tail));

	cby_1__1_ cby_12__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__135_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__7_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__179_ccff_tail),
		.chany_bottom_out(cby_1__1__143_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__143_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__143_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__143_ccff_tail));

	cby_1__1_ cby_13__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__8_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__136_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__180_ccff_tail),
		.chany_bottom_out(cby_1__1__144_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__144_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__144_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__144_ccff_tail));

	cby_1__1_ cby_13__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__136_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__137_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__181_ccff_tail),
		.chany_bottom_out(cby_1__1__145_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__145_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__145_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__145_ccff_tail));

	cby_1__1_ cby_13__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__137_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__138_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__182_ccff_tail),
		.chany_bottom_out(cby_1__1__146_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__146_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__146_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__146_ccff_tail));

	cby_1__1_ cby_13__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__138_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__139_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__183_ccff_tail),
		.chany_bottom_out(cby_1__1__147_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__147_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__147_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__147_ccff_tail));

	cby_1__1_ cby_13__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__139_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__140_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__184_ccff_tail),
		.chany_bottom_out(cby_1__1__148_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__148_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__148_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__148_ccff_tail));

	cby_1__1_ cby_13__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__140_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__141_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__185_ccff_tail),
		.chany_bottom_out(cby_1__1__149_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__149_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__149_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__149_ccff_tail));

	cby_1__1_ cby_13__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__141_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__142_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__186_ccff_tail),
		.chany_bottom_out(cby_1__1__150_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__150_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__150_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__150_ccff_tail));

	cby_1__1_ cby_13__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__142_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__143_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__187_ccff_tail),
		.chany_bottom_out(cby_1__1__151_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__151_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__151_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__151_ccff_tail));

	cby_1__1_ cby_13__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__143_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__144_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__188_ccff_tail),
		.chany_bottom_out(cby_1__1__152_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__152_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__152_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__152_ccff_tail));

	cby_1__1_ cby_13__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__144_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__145_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__189_ccff_tail),
		.chany_bottom_out(cby_1__1__153_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__153_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__153_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__153_ccff_tail));

	cby_1__1_ cby_13__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__145_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__146_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__190_ccff_tail),
		.chany_bottom_out(cby_1__1__154_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__154_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__154_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__154_ccff_tail));

	cby_1__1_ cby_13__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__146_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__147_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__191_ccff_tail),
		.chany_bottom_out(cby_1__1__155_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__155_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__155_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__155_ccff_tail));

	cby_1__1_ cby_13__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__147_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__148_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__192_ccff_tail),
		.chany_bottom_out(cby_1__1__156_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__156_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__156_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__156_ccff_tail));

	cby_1__1_ cby_13__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__148_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__149_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__193_ccff_tail),
		.chany_bottom_out(cby_1__1__157_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__157_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__157_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__157_ccff_tail));

	cby_1__1_ cby_13__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__149_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__150_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__194_ccff_tail),
		.chany_bottom_out(cby_1__1__158_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__158_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__158_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__158_ccff_tail));

	cby_1__1_ cby_13__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__150_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__151_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__195_ccff_tail),
		.chany_bottom_out(cby_1__1__159_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__159_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__159_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__159_ccff_tail));

	cby_1__1_ cby_13__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__151_chany_top_out[0:63]),
		.chany_top_in(sb_1__1__152_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__196_ccff_tail),
		.chany_bottom_out(cby_1__1__160_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__160_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__160_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__160_ccff_tail));

	cby_1__1_ cby_13__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__152_chany_top_out[0:63]),
		.chany_top_in(sb_1__18__8_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__197_ccff_tail),
		.chany_bottom_out(cby_1__1__161_chany_bottom_out[0:63]),
		.chany_top_out(cby_1__1__161_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__161_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_1__1__161_ccff_tail));

	cby_3__1_ cby_3__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__0__0_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__36_ccff_tail),
		.chany_bottom_out(cby_3__1__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__0_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__0_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__0_ccff_tail));

	cby_3__1_ cby_3__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__1_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__2_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__38_ccff_tail),
		.chany_bottom_out(cby_3__1__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__1_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__1_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__1_ccff_tail));

	cby_3__1_ cby_3__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__3_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__4_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__40_ccff_tail),
		.chany_bottom_out(cby_3__1__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__2_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__2_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__2_ccff_tail));

	cby_3__1_ cby_3__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__5_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__6_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__42_ccff_tail),
		.chany_bottom_out(cby_3__1__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__3_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__3_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__3_ccff_tail));

	cby_3__1_ cby_3__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__7_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__8_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__44_ccff_tail),
		.chany_bottom_out(cby_3__1__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__4_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__4_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__4_ccff_tail));

	cby_3__1_ cby_3__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__9_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__10_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__46_ccff_tail),
		.chany_bottom_out(cby_3__1__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__5_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__5_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__5_ccff_tail));

	cby_3__1_ cby_3__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__11_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__12_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__48_ccff_tail),
		.chany_bottom_out(cby_3__1__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__6_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__6_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__6_ccff_tail));

	cby_3__1_ cby_3__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__13_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__14_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__50_ccff_tail),
		.chany_bottom_out(cby_3__1__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__7_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__7_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__7_ccff_tail));

	cby_3__1_ cby_3__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__15_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__16_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__52_ccff_tail),
		.chany_bottom_out(cby_3__1__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__8_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__8_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__8_ccff_tail));

	cby_3__1_ cby_10__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__0__1_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__17_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__144_ccff_tail),
		.chany_bottom_out(cby_3__1__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__9_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__9_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__9_ccff_tail));

	cby_3__1_ cby_10__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__18_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__19_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__146_ccff_tail),
		.chany_bottom_out(cby_3__1__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__10_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__10_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__10_ccff_tail));

	cby_3__1_ cby_10__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__20_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__21_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__148_ccff_tail),
		.chany_bottom_out(cby_3__1__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__11_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__11_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__11_ccff_tail));

	cby_3__1_ cby_10__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__22_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__23_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__150_ccff_tail),
		.chany_bottom_out(cby_3__1__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__12_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__12_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__12_ccff_tail));

	cby_3__1_ cby_10__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__24_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__25_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__152_ccff_tail),
		.chany_bottom_out(cby_3__1__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__13_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__13_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__13_ccff_tail));

	cby_3__1_ cby_10__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__26_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__27_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__154_ccff_tail),
		.chany_bottom_out(cby_3__1__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__14_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__14_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__14_ccff_tail));

	cby_3__1_ cby_10__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__28_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__29_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__156_ccff_tail),
		.chany_bottom_out(cby_3__1__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__15_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__15_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__15_ccff_tail));

	cby_3__1_ cby_10__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__30_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__31_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__158_ccff_tail),
		.chany_bottom_out(cby_3__1__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__16_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__16_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__16_ccff_tail));

	cby_3__1_ cby_10__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__32_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__33_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__160_ccff_tail),
		.chany_bottom_out(cby_3__1__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__1__17_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_waddr_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_raddr_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_(cby_3__1__17_right_grid_left_width_0_height_0_subtile_0__pin_data_in_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__1__17_ccff_tail));

	cby_3__2_ cby_3__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__0_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__37_ccff_tail),
		.chany_bottom_out(cby_3__2__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__0_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__0_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__0_ccff_tail));

	cby_3__2_ cby_3__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__2_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__3_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__39_ccff_tail),
		.chany_bottom_out(cby_3__2__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__1_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__1_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__1_ccff_tail));

	cby_3__2_ cby_3__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__4_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__5_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__41_ccff_tail),
		.chany_bottom_out(cby_3__2__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__2_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__2_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__2_ccff_tail));

	cby_3__2_ cby_3__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__6_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__7_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__43_ccff_tail),
		.chany_bottom_out(cby_3__2__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__3_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__3_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__3_ccff_tail));

	cby_3__2_ cby_3__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__8_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__9_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__45_ccff_tail),
		.chany_bottom_out(cby_3__2__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__4_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__4_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__4_ccff_tail));

	cby_3__2_ cby_3__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__10_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__11_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__47_ccff_tail),
		.chany_bottom_out(cby_3__2__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__5_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__5_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__5_ccff_tail));

	cby_3__2_ cby_3__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__12_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__13_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__49_ccff_tail),
		.chany_bottom_out(cby_3__2__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__6_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__6_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__6_ccff_tail));

	cby_3__2_ cby_3__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__14_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__15_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__51_ccff_tail),
		.chany_bottom_out(cby_3__2__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__7_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__7_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__7_ccff_tail));

	cby_3__2_ cby_3__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__16_chany_top_out[0:63]),
		.chany_top_in(sb_3__18__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__53_ccff_tail),
		.chany_bottom_out(cby_3__2__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__8_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__8_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__8_ccff_tail));

	cby_3__2_ cby_10__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__17_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__18_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__145_ccff_tail),
		.chany_bottom_out(cby_3__2__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__9_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__9_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__9_ccff_tail));

	cby_3__2_ cby_10__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__19_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__20_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__147_ccff_tail),
		.chany_bottom_out(cby_3__2__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__10_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__10_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__10_ccff_tail));

	cby_3__2_ cby_10__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__21_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__22_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__149_ccff_tail),
		.chany_bottom_out(cby_3__2__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__11_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__11_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__11_ccff_tail));

	cby_3__2_ cby_10__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__23_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__24_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__151_ccff_tail),
		.chany_bottom_out(cby_3__2__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__12_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__12_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__12_ccff_tail));

	cby_3__2_ cby_10__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__25_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__26_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__153_ccff_tail),
		.chany_bottom_out(cby_3__2__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__13_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__13_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__13_ccff_tail));

	cby_3__2_ cby_10__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__27_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__28_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__155_ccff_tail),
		.chany_bottom_out(cby_3__2__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__14_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__14_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__14_ccff_tail));

	cby_3__2_ cby_10__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__29_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__30_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__157_ccff_tail),
		.chany_bottom_out(cby_3__2__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__15_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__15_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__15_ccff_tail));

	cby_3__2_ cby_10__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__31_chany_top_out[0:63]),
		.chany_top_in(sb_3__1__32_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__159_ccff_tail),
		.chany_bottom_out(cby_3__2__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__16_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__16_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__16_ccff_tail));

	cby_3__2_ cby_10__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__33_chany_top_out[0:63]),
		.chany_top_in(sb_3__18__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__161_ccff_tail),
		.chany_bottom_out(cby_3__2__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_3__2__17_chany_top_out[0:63]),
		.right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_waddr_7_),
		.right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_raddr_6_),
		.right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_(cby_3__2__17_right_grid_left_width_0_height_1_subtile_0__pin_data_in_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_3__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_3__2__17_ccff_tail));

	cby_4__1_ cby_4__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__0__0_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__0__0_ccff_tail),
		.chany_bottom_out(cby_4__1__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__0_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__0_ccff_tail));

	cby_4__1_ cby_4__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__0_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__0_ccff_tail),
		.chany_bottom_out(cby_4__1__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__1_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__1_ccff_tail));

	cby_4__1_ cby_4__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__1_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__2_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__0_ccff_tail),
		.chany_bottom_out(cby_4__1__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__2_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__2_ccff_tail));

	cby_4__1_ cby_4__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__2_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__3_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__1_ccff_tail),
		.chany_bottom_out(cby_4__1__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__3_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__3_ccff_tail));

	cby_4__1_ cby_4__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__3_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__4_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__1_ccff_tail),
		.chany_bottom_out(cby_4__1__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__4_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__4_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__4_ccff_tail));

	cby_4__1_ cby_4__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__4_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__5_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__2_ccff_tail),
		.chany_bottom_out(cby_4__1__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__5_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__5_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__5_ccff_tail));

	cby_4__1_ cby_4__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__5_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__6_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__2_ccff_tail),
		.chany_bottom_out(cby_4__1__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__6_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__6_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__6_ccff_tail));

	cby_4__1_ cby_4__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__6_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__7_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__3_ccff_tail),
		.chany_bottom_out(cby_4__1__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__7_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__7_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__7_ccff_tail));

	cby_4__1_ cby_4__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__7_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__8_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__3_ccff_tail),
		.chany_bottom_out(cby_4__1__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__8_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__8_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__8_ccff_tail));

	cby_4__1_ cby_4__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__8_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__9_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__4_ccff_tail),
		.chany_bottom_out(cby_4__1__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__9_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__9_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__9_ccff_tail));

	cby_4__1_ cby_4__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__9_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__10_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__4_ccff_tail),
		.chany_bottom_out(cby_4__1__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__10_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__10_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__10_ccff_tail));

	cby_4__1_ cby_4__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__10_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__11_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__5_ccff_tail),
		.chany_bottom_out(cby_4__1__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__11_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__11_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__11_ccff_tail));

	cby_4__1_ cby_4__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__11_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__12_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__5_ccff_tail),
		.chany_bottom_out(cby_4__1__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__12_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__12_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__12_ccff_tail));

	cby_4__1_ cby_4__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__12_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__13_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__6_ccff_tail),
		.chany_bottom_out(cby_4__1__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__13_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__13_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__13_ccff_tail));

	cby_4__1_ cby_4__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__13_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__14_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__6_ccff_tail),
		.chany_bottom_out(cby_4__1__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__14_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__14_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__14_ccff_tail));

	cby_4__1_ cby_4__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__14_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__15_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__7_ccff_tail),
		.chany_bottom_out(cby_4__1__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__15_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__15_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__15_ccff_tail));

	cby_4__1_ cby_4__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__15_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__16_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__7_ccff_tail),
		.chany_bottom_out(cby_4__1__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__16_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__16_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__16_ccff_tail));

	cby_4__1_ cby_4__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__16_chany_top_out[0:63]),
		.chany_top_in(sb_4__18__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__8_ccff_tail),
		.chany_bottom_out(cby_4__1__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__17_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__17_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__17_ccff_tail));

	cby_4__1_ cby_11__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__0__1_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__17_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__0__1_ccff_tail),
		.chany_bottom_out(cby_4__1__18_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__18_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__18_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__18_ccff_tail));

	cby_4__1_ cby_11__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__17_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__18_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__9_ccff_tail),
		.chany_bottom_out(cby_4__1__19_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__19_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__19_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__19_ccff_tail));

	cby_4__1_ cby_11__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__18_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__19_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__8_ccff_tail),
		.chany_bottom_out(cby_4__1__20_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__20_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__20_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__20_ccff_tail));

	cby_4__1_ cby_11__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__19_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__20_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__10_ccff_tail),
		.chany_bottom_out(cby_4__1__21_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__21_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__21_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__21_ccff_tail));

	cby_4__1_ cby_11__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__20_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__21_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__9_ccff_tail),
		.chany_bottom_out(cby_4__1__22_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__22_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__22_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__22_ccff_tail));

	cby_4__1_ cby_11__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__21_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__22_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__11_ccff_tail),
		.chany_bottom_out(cby_4__1__23_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__23_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__23_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__23_ccff_tail));

	cby_4__1_ cby_11__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__22_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__23_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__10_ccff_tail),
		.chany_bottom_out(cby_4__1__24_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__24_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__24_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__24_ccff_tail));

	cby_4__1_ cby_11__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__23_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__24_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__12_ccff_tail),
		.chany_bottom_out(cby_4__1__25_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__25_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__25_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__25_ccff_tail));

	cby_4__1_ cby_11__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__24_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__25_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__11_ccff_tail),
		.chany_bottom_out(cby_4__1__26_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__26_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__26_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__26_ccff_tail));

	cby_4__1_ cby_11__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__25_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__26_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__13_ccff_tail),
		.chany_bottom_out(cby_4__1__27_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__27_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__27_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__27_ccff_tail));

	cby_4__1_ cby_11__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__26_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__27_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__12_ccff_tail),
		.chany_bottom_out(cby_4__1__28_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__28_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__28_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__28_ccff_tail));

	cby_4__1_ cby_11__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__27_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__28_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__14_ccff_tail),
		.chany_bottom_out(cby_4__1__29_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__29_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__29_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__29_ccff_tail));

	cby_4__1_ cby_11__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__28_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__29_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__13_ccff_tail),
		.chany_bottom_out(cby_4__1__30_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__30_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__30_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(ccff_tail[8]));

	cby_4__1_ cby_11__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__29_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__30_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__15_ccff_tail),
		.chany_bottom_out(cby_4__1__31_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__31_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__31_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__31_ccff_tail));

	cby_4__1_ cby_11__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__30_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__31_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__14_ccff_tail),
		.chany_bottom_out(cby_4__1__32_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__32_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__32_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__32_ccff_tail));

	cby_4__1_ cby_11__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__31_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__32_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__16_ccff_tail),
		.chany_bottom_out(cby_4__1__33_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__33_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__33_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__33_ccff_tail));

	cby_4__1_ cby_11__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__32_chany_top_out[0:63]),
		.chany_top_in(sb_4__1__33_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__2__15_ccff_tail),
		.chany_bottom_out(cby_4__1__34_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__34_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__34_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__34_ccff_tail));

	cby_4__1_ cby_11__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__33_chany_top_out[0:63]),
		.chany_top_in(sb_4__18__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_4__1__17_ccff_tail),
		.chany_bottom_out(cby_4__1__35_chany_bottom_out[0:63]),
		.chany_top_out(cby_4__1__35_chany_top_out[0:63]),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_4__1__35_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_4__1__35_ccff_tail));

	cby_14__1_ cby_14__1_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__0__0_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__198_ccff_tail),
		.chany_bottom_out(cby_14__1__0_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__0_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(ccff_tail[1]));

	cby_14__1_ cby_14__2_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__0_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__1_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__199_ccff_tail),
		.chany_bottom_out(cby_14__1__1_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__1_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__1_ccff_tail));

	cby_14__1_ cby_14__3_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__1_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__2_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__200_ccff_tail),
		.chany_bottom_out(cby_14__1__2_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__2_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__2_ccff_tail));

	cby_14__1_ cby_14__4_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__2_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__3_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__201_ccff_tail),
		.chany_bottom_out(cby_14__1__3_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__3_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__3_ccff_tail));

	cby_14__1_ cby_14__5_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__3_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__4_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__202_ccff_tail),
		.chany_bottom_out(cby_14__1__4_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__4_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__4_ccff_tail));

	cby_14__1_ cby_14__6_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__4_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__5_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__203_ccff_tail),
		.chany_bottom_out(cby_14__1__5_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__5_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__5_ccff_tail));

	cby_14__1_ cby_14__7_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__5_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__6_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__204_ccff_tail),
		.chany_bottom_out(cby_14__1__6_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__6_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__6_ccff_tail));

	cby_14__1_ cby_14__8_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__6_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__7_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__205_ccff_tail),
		.chany_bottom_out(cby_14__1__7_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__7_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__7_ccff_tail));

	cby_14__1_ cby_14__9_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__7_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__8_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__206_ccff_tail),
		.chany_bottom_out(cby_14__1__8_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__8_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__8_ccff_tail));

	cby_14__1_ cby_14__10_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__8_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__9_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__207_ccff_tail),
		.chany_bottom_out(cby_14__1__9_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__9_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__9_ccff_tail));

	cby_14__1_ cby_14__11_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__9_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__10_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__208_ccff_tail),
		.chany_bottom_out(cby_14__1__10_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__10_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__10_ccff_tail));

	cby_14__1_ cby_14__12_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__10_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__11_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__209_ccff_tail),
		.chany_bottom_out(cby_14__1__11_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__11_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__11_ccff_tail));

	cby_14__1_ cby_14__13_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__11_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__12_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__210_ccff_tail),
		.chany_bottom_out(cby_14__1__12_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__12_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__12_ccff_tail));

	cby_14__1_ cby_14__14_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__12_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__13_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__211_ccff_tail),
		.chany_bottom_out(cby_14__1__13_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__13_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__13_ccff_tail));

	cby_14__1_ cby_14__15_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__13_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__14_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__212_ccff_tail),
		.chany_bottom_out(cby_14__1__14_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__14_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__14_ccff_tail));

	cby_14__1_ cby_14__16_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__14_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__15_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__213_ccff_tail),
		.chany_bottom_out(cby_14__1__15_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__15_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__15_ccff_tail));

	cby_14__1_ cby_14__17_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__15_chany_top_out[0:63]),
		.chany_top_in(sb_14__1__16_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__214_ccff_tail),
		.chany_bottom_out(cby_14__1__16_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__16_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__16_ccff_tail));

	cby_14__1_ cby_14__18_ (
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_14__1__16_chany_top_out[0:63]),
		.chany_top_in(sb_14__18__0_chany_bottom_out[0:63]),
		.ccff_head(cbx_1__0__215_ccff_tail),
		.chany_bottom_out(cby_14__1__17_chany_bottom_out[0:63]),
		.chany_top_out(cby_14__1__17_chany_top_out[0:63]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_14__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_14__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.ccff_tail(cby_14__1__17_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_29_out));

	direct_interc direct_interc_30_ (
		.in(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_30_out));

	direct_interc direct_interc_31_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_31_out));

	direct_interc direct_interc_32_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_32_out));

	direct_interc direct_interc_33_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_33_out));

	direct_interc direct_interc_34_ (
		.in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_34_out));

	direct_interc direct_interc_35_ (
		.in(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_35_out));

	direct_interc direct_interc_36_ (
		.in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_36_out));

	direct_interc direct_interc_37_ (
		.in(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_37_out));

	direct_interc direct_interc_38_ (
		.in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_38_out));

	direct_interc direct_interc_39_ (
		.in(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_39_out));

	direct_interc direct_interc_40_ (
		.in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_40_out));

	direct_interc direct_interc_41_ (
		.in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_41_out));

	direct_interc direct_interc_42_ (
		.in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_42_out));

	direct_interc direct_interc_43_ (
		.in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_43_out));

	direct_interc direct_interc_44_ (
		.in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_44_out));

	direct_interc direct_interc_45_ (
		.in(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_45_out));

	direct_interc direct_interc_46_ (
		.in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_46_out));

	direct_interc direct_interc_47_ (
		.in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_47_out));

	direct_interc direct_interc_48_ (
		.in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_48_out));

	direct_interc direct_interc_49_ (
		.in(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_49_out));

	direct_interc direct_interc_50_ (
		.in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_50_out));

	direct_interc direct_interc_51_ (
		.in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_51_out));

	direct_interc direct_interc_52_ (
		.in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_52_out));

	direct_interc direct_interc_53_ (
		.in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_53_out));

	direct_interc direct_interc_54_ (
		.in(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_54_out));

	direct_interc direct_interc_55_ (
		.in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_55_out));

	direct_interc direct_interc_56_ (
		.in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_56_out));

	direct_interc direct_interc_57_ (
		.in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_57_out));

	direct_interc direct_interc_58_ (
		.in(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_58_out));

	direct_interc direct_interc_59_ (
		.in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_59_out));

	direct_interc direct_interc_60_ (
		.in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_60_out));

	direct_interc direct_interc_61_ (
		.in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_61_out));

	direct_interc direct_interc_62_ (
		.in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_62_out));

	direct_interc direct_interc_63_ (
		.in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_63_out));

	direct_interc direct_interc_64_ (
		.in(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_64_out));

	direct_interc direct_interc_65_ (
		.in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_65_out));

	direct_interc direct_interc_66_ (
		.in(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_66_out));

	direct_interc direct_interc_67_ (
		.in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_67_out));

	direct_interc direct_interc_68_ (
		.in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_68_out));

	direct_interc direct_interc_69_ (
		.in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_69_out));

	direct_interc direct_interc_70_ (
		.in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_70_out));

	direct_interc direct_interc_71_ (
		.in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_71_out));

	direct_interc direct_interc_72_ (
		.in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_72_out));

	direct_interc direct_interc_73_ (
		.in(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_73_out));

	direct_interc direct_interc_74_ (
		.in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_74_out));

	direct_interc direct_interc_75_ (
		.in(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_75_out));

	direct_interc direct_interc_76_ (
		.in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_76_out));

	direct_interc direct_interc_77_ (
		.in(grid_clb_82_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_77_out));

	direct_interc direct_interc_78_ (
		.in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_78_out));

	direct_interc direct_interc_79_ (
		.in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_79_out));

	direct_interc direct_interc_80_ (
		.in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_80_out));

	direct_interc direct_interc_81_ (
		.in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_81_out));

	direct_interc direct_interc_82_ (
		.in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_82_out));

	direct_interc direct_interc_83_ (
		.in(grid_clb_88_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_83_out));

	direct_interc direct_interc_84_ (
		.in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_84_out));

	direct_interc direct_interc_85_ (
		.in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_85_out));

	direct_interc direct_interc_86_ (
		.in(grid_clb_92_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_86_out));

	direct_interc direct_interc_87_ (
		.in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_87_out));

	direct_interc direct_interc_88_ (
		.in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_88_out));

	direct_interc direct_interc_89_ (
		.in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_89_out));

	direct_interc direct_interc_90_ (
		.in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_90_out));

	direct_interc direct_interc_91_ (
		.in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_91_out));

	direct_interc direct_interc_92_ (
		.in(grid_clb_98_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_92_out));

	direct_interc direct_interc_93_ (
		.in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_93_out));

	direct_interc direct_interc_94_ (
		.in(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_94_out));

	direct_interc direct_interc_95_ (
		.in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_95_out));

	direct_interc direct_interc_96_ (
		.in(grid_clb_102_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_96_out));

	direct_interc direct_interc_97_ (
		.in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_97_out));

	direct_interc direct_interc_98_ (
		.in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_98_out));

	direct_interc direct_interc_99_ (
		.in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_99_out));

	direct_interc direct_interc_100_ (
		.in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_100_out));

	direct_interc direct_interc_101_ (
		.in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_101_out));

	direct_interc direct_interc_102_ (
		.in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_102_out));

	direct_interc direct_interc_103_ (
		.in(grid_clb_110_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_103_out));

	direct_interc direct_interc_104_ (
		.in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_104_out));

	direct_interc direct_interc_105_ (
		.in(grid_clb_112_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_105_out));

	direct_interc direct_interc_106_ (
		.in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_106_out));

	direct_interc direct_interc_107_ (
		.in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_107_out));

	direct_interc direct_interc_108_ (
		.in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_108_out));

	direct_interc direct_interc_109_ (
		.in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_109_out));

	direct_interc direct_interc_110_ (
		.in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_110_out));

	direct_interc direct_interc_111_ (
		.in(grid_clb_118_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_111_out));

	direct_interc direct_interc_112_ (
		.in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_112_out));

	direct_interc direct_interc_113_ (
		.in(grid_clb_120_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_113_out));

	direct_interc direct_interc_114_ (
		.in(grid_clb_121_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_114_out));

	direct_interc direct_interc_115_ (
		.in(grid_clb_122_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_115_out));

	direct_interc direct_interc_116_ (
		.in(grid_clb_123_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_116_out));

	direct_interc direct_interc_117_ (
		.in(grid_clb_124_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_117_out));

	direct_interc direct_interc_118_ (
		.in(grid_clb_125_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_118_out));

	direct_interc direct_interc_119_ (
		.in(grid_clb_127_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_119_out));

	direct_interc direct_interc_120_ (
		.in(grid_clb_128_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_120_out));

	direct_interc direct_interc_121_ (
		.in(grid_clb_129_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_121_out));

	direct_interc direct_interc_122_ (
		.in(grid_clb_130_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_122_out));

	direct_interc direct_interc_123_ (
		.in(grid_clb_131_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_123_out));

	direct_interc direct_interc_124_ (
		.in(grid_clb_132_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_124_out));

	direct_interc direct_interc_125_ (
		.in(grid_clb_133_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_125_out));

	direct_interc direct_interc_126_ (
		.in(grid_clb_134_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_126_out));

	direct_interc direct_interc_127_ (
		.in(grid_clb_135_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_127_out));

	direct_interc direct_interc_128_ (
		.in(grid_clb_136_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_128_out));

	direct_interc direct_interc_129_ (
		.in(grid_clb_137_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_129_out));

	direct_interc direct_interc_130_ (
		.in(grid_clb_138_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_130_out));

	direct_interc direct_interc_131_ (
		.in(grid_clb_139_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_131_out));

	direct_interc direct_interc_132_ (
		.in(grid_clb_140_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_132_out));

	direct_interc direct_interc_133_ (
		.in(grid_clb_141_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_133_out));

	direct_interc direct_interc_134_ (
		.in(grid_clb_142_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_134_out));

	direct_interc direct_interc_135_ (
		.in(grid_clb_143_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_135_out));

	direct_interc direct_interc_136_ (
		.in(grid_clb_145_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_136_out));

	direct_interc direct_interc_137_ (
		.in(grid_clb_146_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_137_out));

	direct_interc direct_interc_138_ (
		.in(grid_clb_147_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_138_out));

	direct_interc direct_interc_139_ (
		.in(grid_clb_148_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_139_out));

	direct_interc direct_interc_140_ (
		.in(grid_clb_149_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_140_out));

	direct_interc direct_interc_141_ (
		.in(grid_clb_150_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_141_out));

	direct_interc direct_interc_142_ (
		.in(grid_clb_151_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_142_out));

	direct_interc direct_interc_143_ (
		.in(grid_clb_152_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_143_out));

	direct_interc direct_interc_144_ (
		.in(grid_clb_153_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_144_out));

	direct_interc direct_interc_145_ (
		.in(grid_clb_154_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_145_out));

	direct_interc direct_interc_146_ (
		.in(grid_clb_155_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_146_out));

	direct_interc direct_interc_147_ (
		.in(grid_clb_156_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_147_out));

	direct_interc direct_interc_148_ (
		.in(grid_clb_157_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_148_out));

	direct_interc direct_interc_149_ (
		.in(grid_clb_158_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_149_out));

	direct_interc direct_interc_150_ (
		.in(grid_clb_159_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_150_out));

	direct_interc direct_interc_151_ (
		.in(grid_clb_160_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_151_out));

	direct_interc direct_interc_152_ (
		.in(grid_clb_161_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_152_out));

	direct_interc direct_interc_153_ (
		.in(grid_clb_163_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_153_out));

	direct_interc direct_interc_154_ (
		.in(grid_clb_164_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_154_out));

	direct_interc direct_interc_155_ (
		.in(grid_clb_165_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_155_out));

	direct_interc direct_interc_156_ (
		.in(grid_clb_166_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_156_out));

	direct_interc direct_interc_157_ (
		.in(grid_clb_167_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_157_out));

	direct_interc direct_interc_158_ (
		.in(grid_clb_168_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_158_out));

	direct_interc direct_interc_159_ (
		.in(grid_clb_169_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_159_out));

	direct_interc direct_interc_160_ (
		.in(grid_clb_170_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_160_out));

	direct_interc direct_interc_161_ (
		.in(grid_clb_171_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_161_out));

	direct_interc direct_interc_162_ (
		.in(grid_clb_172_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_162_out));

	direct_interc direct_interc_163_ (
		.in(grid_clb_173_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_163_out));

	direct_interc direct_interc_164_ (
		.in(grid_clb_174_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_164_out));

	direct_interc direct_interc_165_ (
		.in(grid_clb_175_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_165_out));

	direct_interc direct_interc_166_ (
		.in(grid_clb_176_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_166_out));

	direct_interc direct_interc_167_ (
		.in(grid_clb_177_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_167_out));

	direct_interc direct_interc_168_ (
		.in(grid_clb_178_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_168_out));

	direct_interc direct_interc_169_ (
		.in(grid_clb_179_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_169_out));

	direct_interc direct_interc_170_ (
		.in(grid_clb_181_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_170_out));

	direct_interc direct_interc_171_ (
		.in(grid_clb_182_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_171_out));

	direct_interc direct_interc_172_ (
		.in(grid_clb_183_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_172_out));

	direct_interc direct_interc_173_ (
		.in(grid_clb_184_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_173_out));

	direct_interc direct_interc_174_ (
		.in(grid_clb_185_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_174_out));

	direct_interc direct_interc_175_ (
		.in(grid_clb_186_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_175_out));

	direct_interc direct_interc_176_ (
		.in(grid_clb_187_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_176_out));

	direct_interc direct_interc_177_ (
		.in(grid_clb_188_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_177_out));

	direct_interc direct_interc_178_ (
		.in(grid_clb_189_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_178_out));

	direct_interc direct_interc_179_ (
		.in(grid_clb_190_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_179_out));

	direct_interc direct_interc_180_ (
		.in(grid_clb_191_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_180_out));

	direct_interc direct_interc_181_ (
		.in(grid_clb_192_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_181_out));

	direct_interc direct_interc_182_ (
		.in(grid_clb_193_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_182_out));

	direct_interc direct_interc_183_ (
		.in(grid_clb_194_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_183_out));

	direct_interc direct_interc_184_ (
		.in(grid_clb_195_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_184_out));

	direct_interc direct_interc_185_ (
		.in(grid_clb_196_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_185_out));

	direct_interc direct_interc_186_ (
		.in(grid_clb_197_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_186_out));

	direct_interc direct_interc_187_ (
		.in(grid_clb_199_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_187_out));

	direct_interc direct_interc_188_ (
		.in(grid_clb_200_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_188_out));

	direct_interc direct_interc_189_ (
		.in(grid_clb_201_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_189_out));

	direct_interc direct_interc_190_ (
		.in(grid_clb_202_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_190_out));

	direct_interc direct_interc_191_ (
		.in(grid_clb_203_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_191_out));

	direct_interc direct_interc_192_ (
		.in(grid_clb_204_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_192_out));

	direct_interc direct_interc_193_ (
		.in(grid_clb_205_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_193_out));

	direct_interc direct_interc_194_ (
		.in(grid_clb_206_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_194_out));

	direct_interc direct_interc_195_ (
		.in(grid_clb_207_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_195_out));

	direct_interc direct_interc_196_ (
		.in(grid_clb_208_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_196_out));

	direct_interc direct_interc_197_ (
		.in(grid_clb_209_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_197_out));

	direct_interc direct_interc_198_ (
		.in(grid_clb_210_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_198_out));

	direct_interc direct_interc_199_ (
		.in(grid_clb_211_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_199_out));

	direct_interc direct_interc_200_ (
		.in(grid_clb_212_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_200_out));

	direct_interc direct_interc_201_ (
		.in(grid_clb_213_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_201_out));

	direct_interc direct_interc_202_ (
		.in(grid_clb_214_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_202_out));

	direct_interc direct_interc_203_ (
		.in(grid_clb_215_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_203_out));

	direct_interc direct_interc_204_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_204_out));

	direct_interc direct_interc_205_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_205_out));

	direct_interc direct_interc_206_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_206_out));

	direct_interc direct_interc_207_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_207_out));

	direct_interc direct_interc_208_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_208_out));

	direct_interc direct_interc_209_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_209_out));

	direct_interc direct_interc_210_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_210_out));

	direct_interc direct_interc_211_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_211_out));

	direct_interc direct_interc_212_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_212_out));

	direct_interc direct_interc_213_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_213_out));

	direct_interc direct_interc_214_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_214_out));

	direct_interc direct_interc_215_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_215_out));

	direct_interc direct_interc_216_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_216_out));

	direct_interc direct_interc_217_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_217_out));

	direct_interc direct_interc_218_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_218_out));

	direct_interc direct_interc_219_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_219_out));

	direct_interc direct_interc_220_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_220_out));

	direct_interc direct_interc_221_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_221_out));

	direct_interc direct_interc_222_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_222_out));

	direct_interc direct_interc_223_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_223_out));

	direct_interc direct_interc_224_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_224_out));

	direct_interc direct_interc_225_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_225_out));

	direct_interc direct_interc_226_ (
		.in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_226_out));

	direct_interc direct_interc_227_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_227_out));

	direct_interc direct_interc_228_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_228_out));

	direct_interc direct_interc_229_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_229_out));

	direct_interc direct_interc_230_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_230_out));

	direct_interc direct_interc_231_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_231_out));

	direct_interc direct_interc_232_ (
		.in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_232_out));

	direct_interc direct_interc_233_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_233_out));

	direct_interc direct_interc_234_ (
		.in(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_234_out));

	direct_interc direct_interc_235_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_235_out));

	direct_interc direct_interc_236_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_236_out));

	direct_interc direct_interc_237_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_237_out));

	direct_interc direct_interc_238_ (
		.in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_238_out));

	direct_interc direct_interc_239_ (
		.in(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_239_out));

	direct_interc direct_interc_240_ (
		.in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_240_out));

	direct_interc direct_interc_241_ (
		.in(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_241_out));

	direct_interc direct_interc_242_ (
		.in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_242_out));

	direct_interc direct_interc_243_ (
		.in(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_243_out));

	direct_interc direct_interc_244_ (
		.in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_244_out));

	direct_interc direct_interc_245_ (
		.in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_245_out));

	direct_interc direct_interc_246_ (
		.in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_246_out));

	direct_interc direct_interc_247_ (
		.in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_247_out));

	direct_interc direct_interc_248_ (
		.in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_248_out));

	direct_interc direct_interc_249_ (
		.in(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_249_out));

	direct_interc direct_interc_250_ (
		.in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_250_out));

	direct_interc direct_interc_251_ (
		.in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_251_out));

	direct_interc direct_interc_252_ (
		.in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_252_out));

	direct_interc direct_interc_253_ (
		.in(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_253_out));

	direct_interc direct_interc_254_ (
		.in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_254_out));

	direct_interc direct_interc_255_ (
		.in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_255_out));

	direct_interc direct_interc_256_ (
		.in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_256_out));

	direct_interc direct_interc_257_ (
		.in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_257_out));

	direct_interc direct_interc_258_ (
		.in(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_258_out));

	direct_interc direct_interc_259_ (
		.in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_259_out));

	direct_interc direct_interc_260_ (
		.in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_260_out));

	direct_interc direct_interc_261_ (
		.in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_261_out));

	direct_interc direct_interc_262_ (
		.in(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_262_out));

	direct_interc direct_interc_263_ (
		.in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_263_out));

	direct_interc direct_interc_264_ (
		.in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_264_out));

	direct_interc direct_interc_265_ (
		.in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_265_out));

	direct_interc direct_interc_266_ (
		.in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_266_out));

	direct_interc direct_interc_267_ (
		.in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_267_out));

	direct_interc direct_interc_268_ (
		.in(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_268_out));

	direct_interc direct_interc_269_ (
		.in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_269_out));

	direct_interc direct_interc_270_ (
		.in(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_270_out));

	direct_interc direct_interc_271_ (
		.in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_271_out));

	direct_interc direct_interc_272_ (
		.in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_272_out));

	direct_interc direct_interc_273_ (
		.in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_273_out));

	direct_interc direct_interc_274_ (
		.in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_274_out));

	direct_interc direct_interc_275_ (
		.in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_275_out));

	direct_interc direct_interc_276_ (
		.in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_276_out));

	direct_interc direct_interc_277_ (
		.in(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_277_out));

	direct_interc direct_interc_278_ (
		.in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_278_out));

	direct_interc direct_interc_279_ (
		.in(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_279_out));

	direct_interc direct_interc_280_ (
		.in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_280_out));

	direct_interc direct_interc_281_ (
		.in(grid_clb_82_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_281_out));

	direct_interc direct_interc_282_ (
		.in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_282_out));

	direct_interc direct_interc_283_ (
		.in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_283_out));

	direct_interc direct_interc_284_ (
		.in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_284_out));

	direct_interc direct_interc_285_ (
		.in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_285_out));

	direct_interc direct_interc_286_ (
		.in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_286_out));

	direct_interc direct_interc_287_ (
		.in(grid_clb_88_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_287_out));

	direct_interc direct_interc_288_ (
		.in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_288_out));

	direct_interc direct_interc_289_ (
		.in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_289_out));

	direct_interc direct_interc_290_ (
		.in(grid_clb_92_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_290_out));

	direct_interc direct_interc_291_ (
		.in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_291_out));

	direct_interc direct_interc_292_ (
		.in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_292_out));

	direct_interc direct_interc_293_ (
		.in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_293_out));

	direct_interc direct_interc_294_ (
		.in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_294_out));

	direct_interc direct_interc_295_ (
		.in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_295_out));

	direct_interc direct_interc_296_ (
		.in(grid_clb_98_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_296_out));

	direct_interc direct_interc_297_ (
		.in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_297_out));

	direct_interc direct_interc_298_ (
		.in(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_298_out));

	direct_interc direct_interc_299_ (
		.in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_299_out));

	direct_interc direct_interc_300_ (
		.in(grid_clb_102_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_300_out));

	direct_interc direct_interc_301_ (
		.in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_301_out));

	direct_interc direct_interc_302_ (
		.in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_302_out));

	direct_interc direct_interc_303_ (
		.in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_303_out));

	direct_interc direct_interc_304_ (
		.in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_304_out));

	direct_interc direct_interc_305_ (
		.in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_305_out));

	direct_interc direct_interc_306_ (
		.in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_306_out));

	direct_interc direct_interc_307_ (
		.in(grid_clb_110_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_307_out));

	direct_interc direct_interc_308_ (
		.in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_308_out));

	direct_interc direct_interc_309_ (
		.in(grid_clb_112_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_309_out));

	direct_interc direct_interc_310_ (
		.in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_310_out));

	direct_interc direct_interc_311_ (
		.in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_311_out));

	direct_interc direct_interc_312_ (
		.in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_312_out));

	direct_interc direct_interc_313_ (
		.in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_313_out));

	direct_interc direct_interc_314_ (
		.in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_314_out));

	direct_interc direct_interc_315_ (
		.in(grid_clb_118_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_315_out));

	direct_interc direct_interc_316_ (
		.in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_316_out));

	direct_interc direct_interc_317_ (
		.in(grid_clb_120_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_317_out));

	direct_interc direct_interc_318_ (
		.in(grid_clb_121_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_318_out));

	direct_interc direct_interc_319_ (
		.in(grid_clb_122_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_319_out));

	direct_interc direct_interc_320_ (
		.in(grid_clb_123_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_320_out));

	direct_interc direct_interc_321_ (
		.in(grid_clb_124_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_321_out));

	direct_interc direct_interc_322_ (
		.in(grid_clb_125_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_322_out));

	direct_interc direct_interc_323_ (
		.in(grid_clb_127_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_323_out));

	direct_interc direct_interc_324_ (
		.in(grid_clb_128_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_324_out));

	direct_interc direct_interc_325_ (
		.in(grid_clb_129_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_325_out));

	direct_interc direct_interc_326_ (
		.in(grid_clb_130_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_326_out));

	direct_interc direct_interc_327_ (
		.in(grid_clb_131_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_327_out));

	direct_interc direct_interc_328_ (
		.in(grid_clb_132_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_328_out));

	direct_interc direct_interc_329_ (
		.in(grid_clb_133_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_329_out));

	direct_interc direct_interc_330_ (
		.in(grid_clb_134_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_330_out));

	direct_interc direct_interc_331_ (
		.in(grid_clb_135_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_331_out));

	direct_interc direct_interc_332_ (
		.in(grid_clb_136_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_332_out));

	direct_interc direct_interc_333_ (
		.in(grid_clb_137_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_333_out));

	direct_interc direct_interc_334_ (
		.in(grid_clb_138_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_334_out));

	direct_interc direct_interc_335_ (
		.in(grid_clb_139_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_335_out));

	direct_interc direct_interc_336_ (
		.in(grid_clb_140_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_336_out));

	direct_interc direct_interc_337_ (
		.in(grid_clb_141_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_337_out));

	direct_interc direct_interc_338_ (
		.in(grid_clb_142_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_338_out));

	direct_interc direct_interc_339_ (
		.in(grid_clb_143_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_339_out));

	direct_interc direct_interc_340_ (
		.in(grid_clb_145_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_340_out));

	direct_interc direct_interc_341_ (
		.in(grid_clb_146_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_341_out));

	direct_interc direct_interc_342_ (
		.in(grid_clb_147_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_342_out));

	direct_interc direct_interc_343_ (
		.in(grid_clb_148_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_343_out));

	direct_interc direct_interc_344_ (
		.in(grid_clb_149_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_344_out));

	direct_interc direct_interc_345_ (
		.in(grid_clb_150_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_345_out));

	direct_interc direct_interc_346_ (
		.in(grid_clb_151_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_346_out));

	direct_interc direct_interc_347_ (
		.in(grid_clb_152_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_347_out));

	direct_interc direct_interc_348_ (
		.in(grid_clb_153_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_348_out));

	direct_interc direct_interc_349_ (
		.in(grid_clb_154_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_349_out));

	direct_interc direct_interc_350_ (
		.in(grid_clb_155_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_350_out));

	direct_interc direct_interc_351_ (
		.in(grid_clb_156_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_351_out));

	direct_interc direct_interc_352_ (
		.in(grid_clb_157_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_352_out));

	direct_interc direct_interc_353_ (
		.in(grid_clb_158_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_353_out));

	direct_interc direct_interc_354_ (
		.in(grid_clb_159_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_354_out));

	direct_interc direct_interc_355_ (
		.in(grid_clb_160_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_355_out));

	direct_interc direct_interc_356_ (
		.in(grid_clb_161_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_356_out));

	direct_interc direct_interc_357_ (
		.in(grid_clb_163_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_357_out));

	direct_interc direct_interc_358_ (
		.in(grid_clb_164_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_358_out));

	direct_interc direct_interc_359_ (
		.in(grid_clb_165_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_359_out));

	direct_interc direct_interc_360_ (
		.in(grid_clb_166_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_360_out));

	direct_interc direct_interc_361_ (
		.in(grid_clb_167_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_361_out));

	direct_interc direct_interc_362_ (
		.in(grid_clb_168_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_362_out));

	direct_interc direct_interc_363_ (
		.in(grid_clb_169_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_363_out));

	direct_interc direct_interc_364_ (
		.in(grid_clb_170_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_364_out));

	direct_interc direct_interc_365_ (
		.in(grid_clb_171_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_365_out));

	direct_interc direct_interc_366_ (
		.in(grid_clb_172_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_366_out));

	direct_interc direct_interc_367_ (
		.in(grid_clb_173_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_367_out));

	direct_interc direct_interc_368_ (
		.in(grid_clb_174_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_368_out));

	direct_interc direct_interc_369_ (
		.in(grid_clb_175_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_369_out));

	direct_interc direct_interc_370_ (
		.in(grid_clb_176_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_370_out));

	direct_interc direct_interc_371_ (
		.in(grid_clb_177_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_371_out));

	direct_interc direct_interc_372_ (
		.in(grid_clb_178_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_372_out));

	direct_interc direct_interc_373_ (
		.in(grid_clb_179_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_373_out));

	direct_interc direct_interc_374_ (
		.in(grid_clb_181_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_374_out));

	direct_interc direct_interc_375_ (
		.in(grid_clb_182_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_375_out));

	direct_interc direct_interc_376_ (
		.in(grid_clb_183_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_376_out));

	direct_interc direct_interc_377_ (
		.in(grid_clb_184_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_377_out));

	direct_interc direct_interc_378_ (
		.in(grid_clb_185_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_378_out));

	direct_interc direct_interc_379_ (
		.in(grid_clb_186_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_379_out));

	direct_interc direct_interc_380_ (
		.in(grid_clb_187_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_380_out));

	direct_interc direct_interc_381_ (
		.in(grid_clb_188_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_381_out));

	direct_interc direct_interc_382_ (
		.in(grid_clb_189_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_382_out));

	direct_interc direct_interc_383_ (
		.in(grid_clb_190_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_383_out));

	direct_interc direct_interc_384_ (
		.in(grid_clb_191_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_384_out));

	direct_interc direct_interc_385_ (
		.in(grid_clb_192_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_385_out));

	direct_interc direct_interc_386_ (
		.in(grid_clb_193_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_386_out));

	direct_interc direct_interc_387_ (
		.in(grid_clb_194_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_387_out));

	direct_interc direct_interc_388_ (
		.in(grid_clb_195_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_388_out));

	direct_interc direct_interc_389_ (
		.in(grid_clb_196_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_389_out));

	direct_interc direct_interc_390_ (
		.in(grid_clb_197_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_390_out));

	direct_interc direct_interc_391_ (
		.in(grid_clb_199_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_391_out));

	direct_interc direct_interc_392_ (
		.in(grid_clb_200_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_392_out));

	direct_interc direct_interc_393_ (
		.in(grid_clb_201_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_393_out));

	direct_interc direct_interc_394_ (
		.in(grid_clb_202_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_394_out));

	direct_interc direct_interc_395_ (
		.in(grid_clb_203_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_395_out));

	direct_interc direct_interc_396_ (
		.in(grid_clb_204_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_396_out));

	direct_interc direct_interc_397_ (
		.in(grid_clb_205_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_397_out));

	direct_interc direct_interc_398_ (
		.in(grid_clb_206_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_398_out));

	direct_interc direct_interc_399_ (
		.in(grid_clb_207_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_399_out));

	direct_interc direct_interc_400_ (
		.in(grid_clb_208_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_400_out));

	direct_interc direct_interc_401_ (
		.in(grid_clb_209_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_401_out));

	direct_interc direct_interc_402_ (
		.in(grid_clb_210_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_402_out));

	direct_interc direct_interc_403_ (
		.in(grid_clb_211_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_403_out));

	direct_interc direct_interc_404_ (
		.in(grid_clb_212_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_404_out));

	direct_interc direct_interc_405_ (
		.in(grid_clb_213_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_405_out));

	direct_interc direct_interc_406_ (
		.in(grid_clb_214_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_406_out));

	direct_interc direct_interc_407_ (
		.in(grid_clb_215_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_407_out));

	direct_interc direct_interc_408_ (
		.in(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_408_out));

	direct_interc direct_interc_409_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_409_out));

	direct_interc direct_interc_410_ (
		.in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_410_out));

	direct_interc direct_interc_411_ (
		.in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_411_out));

	direct_interc direct_interc_412_ (
		.in(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_412_out));

	direct_interc direct_interc_413_ (
		.in(grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_413_out));

	direct_interc direct_interc_414_ (
		.in(grid_clb_108_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_414_out));

	direct_interc direct_interc_415_ (
		.in(grid_clb_126_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_415_out));

	direct_interc direct_interc_416_ (
		.in(grid_clb_144_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_416_out));

	direct_interc direct_interc_417_ (
		.in(grid_clb_162_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_417_out));

	direct_interc direct_interc_418_ (
		.in(grid_clb_180_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_418_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
// `default_nettype none




