

module fpga_core
( config_enable, pReset, prog_clk, Test_en, IO_ISOL_N, reset, gfpga_pad_sofa_plus_io_SOC_IN, gfpga_pad_sofa_plus_io_SOC_OUT, gfpga_pad_sofa_plus_io_SOC_DIR, ccff_head, ccff_tail, sc_head, sc_tail, clk0 ); 
  input [0:0] config_enable;
  input [0:0] pReset;
  input [0:0] prog_clk;
  input [0:0] Test_en;
  input [0:0] IO_ISOL_N;
  input [0:0] reset;
  input [0:143] gfpga_pad_sofa_plus_io_SOC_IN;
  output [0:143] gfpga_pad_sofa_plus_io_SOC_OUT;
  output [0:143] gfpga_pad_sofa_plus_io_SOC_DIR;
  input [0:11] ccff_head;
  output [0:11] ccff_tail;
  input sc_head;
  output sc_tail;
  input clk0;

  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__0_ccff_tail;
  wire [0:19] cbx_1__0__0_chanx_left_out;
  wire [0:19] cbx_1__0__0_chanx_right_out;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__10_ccff_tail;
  wire [0:19] cbx_1__0__10_chanx_left_out;
  wire [0:19] cbx_1__0__10_chanx_right_out;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__11_ccff_tail;
  wire [0:19] cbx_1__0__11_chanx_left_out;
  wire [0:19] cbx_1__0__11_chanx_right_out;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__1_ccff_tail;
  wire [0:19] cbx_1__0__1_chanx_left_out;
  wire [0:19] cbx_1__0__1_chanx_right_out;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__2_ccff_tail;
  wire [0:19] cbx_1__0__2_chanx_left_out;
  wire [0:19] cbx_1__0__2_chanx_right_out;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__3_ccff_tail;
  wire [0:19] cbx_1__0__3_chanx_left_out;
  wire [0:19] cbx_1__0__3_chanx_right_out;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__4_ccff_tail;
  wire [0:19] cbx_1__0__4_chanx_left_out;
  wire [0:19] cbx_1__0__4_chanx_right_out;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__5_ccff_tail;
  wire [0:19] cbx_1__0__5_chanx_left_out;
  wire [0:19] cbx_1__0__5_chanx_right_out;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__6_ccff_tail;
  wire [0:19] cbx_1__0__6_chanx_left_out;
  wire [0:19] cbx_1__0__6_chanx_right_out;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__7_ccff_tail;
  wire [0:19] cbx_1__0__7_chanx_left_out;
  wire [0:19] cbx_1__0__7_chanx_right_out;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__8_ccff_tail;
  wire [0:19] cbx_1__0__8_chanx_left_out;
  wire [0:19] cbx_1__0__8_chanx_right_out;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
  wire [0:0] cbx_1__0__9_ccff_tail;
  wire [0:19] cbx_1__0__9_chanx_left_out;
  wire [0:19] cbx_1__0__9_chanx_right_out;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__0_ccff_tail;
  wire [0:19] cbx_1__12__0_chanx_left_out;
  wire [0:19] cbx_1__12__0_chanx_right_out;
  wire [0:0] cbx_1__12__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__10_ccff_tail;
  wire [0:19] cbx_1__12__10_chanx_left_out;
  wire [0:19] cbx_1__12__10_chanx_right_out;
  wire [0:0] cbx_1__12__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__11_ccff_tail;
  wire [0:19] cbx_1__12__11_chanx_left_out;
  wire [0:19] cbx_1__12__11_chanx_right_out;
  wire [0:0] cbx_1__12__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__1_ccff_tail;
  wire [0:19] cbx_1__12__1_chanx_left_out;
  wire [0:19] cbx_1__12__1_chanx_right_out;
  wire [0:0] cbx_1__12__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__2_ccff_tail;
  wire [0:19] cbx_1__12__2_chanx_left_out;
  wire [0:19] cbx_1__12__2_chanx_right_out;
  wire [0:0] cbx_1__12__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__3_ccff_tail;
  wire [0:19] cbx_1__12__3_chanx_left_out;
  wire [0:19] cbx_1__12__3_chanx_right_out;
  wire [0:0] cbx_1__12__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__4_ccff_tail;
  wire [0:19] cbx_1__12__4_chanx_left_out;
  wire [0:19] cbx_1__12__4_chanx_right_out;
  wire [0:0] cbx_1__12__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__5_ccff_tail;
  wire [0:19] cbx_1__12__5_chanx_left_out;
  wire [0:19] cbx_1__12__5_chanx_right_out;
  wire [0:0] cbx_1__12__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__6_ccff_tail;
  wire [0:19] cbx_1__12__6_chanx_left_out;
  wire [0:19] cbx_1__12__6_chanx_right_out;
  wire [0:0] cbx_1__12__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__7_ccff_tail;
  wire [0:19] cbx_1__12__7_chanx_left_out;
  wire [0:19] cbx_1__12__7_chanx_right_out;
  wire [0:0] cbx_1__12__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__8_ccff_tail;
  wire [0:19] cbx_1__12__8_chanx_left_out;
  wire [0:19] cbx_1__12__8_chanx_right_out;
  wire [0:0] cbx_1__12__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__12__9_ccff_tail;
  wire [0:19] cbx_1__12__9_chanx_left_out;
  wire [0:19] cbx_1__12__9_chanx_right_out;
  wire [0:0] cbx_1__12__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__0_ccff_tail;
  wire [0:19] cbx_1__1__0_chanx_left_out;
  wire [0:19] cbx_1__1__0_chanx_right_out;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__100_ccff_tail;
  wire [0:19] cbx_1__1__100_chanx_left_out;
  wire [0:19] cbx_1__1__100_chanx_right_out;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__101_ccff_tail;
  wire [0:19] cbx_1__1__101_chanx_left_out;
  wire [0:19] cbx_1__1__101_chanx_right_out;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__102_ccff_tail;
  wire [0:19] cbx_1__1__102_chanx_left_out;
  wire [0:19] cbx_1__1__102_chanx_right_out;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__103_ccff_tail;
  wire [0:19] cbx_1__1__103_chanx_left_out;
  wire [0:19] cbx_1__1__103_chanx_right_out;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__104_ccff_tail;
  wire [0:19] cbx_1__1__104_chanx_left_out;
  wire [0:19] cbx_1__1__104_chanx_right_out;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__105_ccff_tail;
  wire [0:19] cbx_1__1__105_chanx_left_out;
  wire [0:19] cbx_1__1__105_chanx_right_out;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__106_ccff_tail;
  wire [0:19] cbx_1__1__106_chanx_left_out;
  wire [0:19] cbx_1__1__106_chanx_right_out;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__107_ccff_tail;
  wire [0:19] cbx_1__1__107_chanx_left_out;
  wire [0:19] cbx_1__1__107_chanx_right_out;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__10_ccff_tail;
  wire [0:19] cbx_1__1__10_chanx_left_out;
  wire [0:19] cbx_1__1__10_chanx_right_out;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__11_ccff_tail;
  wire [0:19] cbx_1__1__11_chanx_left_out;
  wire [0:19] cbx_1__1__11_chanx_right_out;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__12_ccff_tail;
  wire [0:19] cbx_1__1__12_chanx_left_out;
  wire [0:19] cbx_1__1__12_chanx_right_out;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__13_ccff_tail;
  wire [0:19] cbx_1__1__13_chanx_left_out;
  wire [0:19] cbx_1__1__13_chanx_right_out;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__14_ccff_tail;
  wire [0:19] cbx_1__1__14_chanx_left_out;
  wire [0:19] cbx_1__1__14_chanx_right_out;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__15_ccff_tail;
  wire [0:19] cbx_1__1__15_chanx_left_out;
  wire [0:19] cbx_1__1__15_chanx_right_out;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__16_ccff_tail;
  wire [0:19] cbx_1__1__16_chanx_left_out;
  wire [0:19] cbx_1__1__16_chanx_right_out;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__17_ccff_tail;
  wire [0:19] cbx_1__1__17_chanx_left_out;
  wire [0:19] cbx_1__1__17_chanx_right_out;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__18_ccff_tail;
  wire [0:19] cbx_1__1__18_chanx_left_out;
  wire [0:19] cbx_1__1__18_chanx_right_out;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__19_ccff_tail;
  wire [0:19] cbx_1__1__19_chanx_left_out;
  wire [0:19] cbx_1__1__19_chanx_right_out;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__1_ccff_tail;
  wire [0:19] cbx_1__1__1_chanx_left_out;
  wire [0:19] cbx_1__1__1_chanx_right_out;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__20_ccff_tail;
  wire [0:19] cbx_1__1__20_chanx_left_out;
  wire [0:19] cbx_1__1__20_chanx_right_out;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__21_ccff_tail;
  wire [0:19] cbx_1__1__21_chanx_left_out;
  wire [0:19] cbx_1__1__21_chanx_right_out;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__22_ccff_tail;
  wire [0:19] cbx_1__1__22_chanx_left_out;
  wire [0:19] cbx_1__1__22_chanx_right_out;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__23_ccff_tail;
  wire [0:19] cbx_1__1__23_chanx_left_out;
  wire [0:19] cbx_1__1__23_chanx_right_out;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__24_ccff_tail;
  wire [0:19] cbx_1__1__24_chanx_left_out;
  wire [0:19] cbx_1__1__24_chanx_right_out;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__25_ccff_tail;
  wire [0:19] cbx_1__1__25_chanx_left_out;
  wire [0:19] cbx_1__1__25_chanx_right_out;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__26_ccff_tail;
  wire [0:19] cbx_1__1__26_chanx_left_out;
  wire [0:19] cbx_1__1__26_chanx_right_out;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__27_ccff_tail;
  wire [0:19] cbx_1__1__27_chanx_left_out;
  wire [0:19] cbx_1__1__27_chanx_right_out;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__28_ccff_tail;
  wire [0:19] cbx_1__1__28_chanx_left_out;
  wire [0:19] cbx_1__1__28_chanx_right_out;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__29_ccff_tail;
  wire [0:19] cbx_1__1__29_chanx_left_out;
  wire [0:19] cbx_1__1__29_chanx_right_out;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__2_ccff_tail;
  wire [0:19] cbx_1__1__2_chanx_left_out;
  wire [0:19] cbx_1__1__2_chanx_right_out;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__30_ccff_tail;
  wire [0:19] cbx_1__1__30_chanx_left_out;
  wire [0:19] cbx_1__1__30_chanx_right_out;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__31_ccff_tail;
  wire [0:19] cbx_1__1__31_chanx_left_out;
  wire [0:19] cbx_1__1__31_chanx_right_out;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__32_ccff_tail;
  wire [0:19] cbx_1__1__32_chanx_left_out;
  wire [0:19] cbx_1__1__32_chanx_right_out;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__33_ccff_tail;
  wire [0:19] cbx_1__1__33_chanx_left_out;
  wire [0:19] cbx_1__1__33_chanx_right_out;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__34_ccff_tail;
  wire [0:19] cbx_1__1__34_chanx_left_out;
  wire [0:19] cbx_1__1__34_chanx_right_out;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__35_ccff_tail;
  wire [0:19] cbx_1__1__35_chanx_left_out;
  wire [0:19] cbx_1__1__35_chanx_right_out;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__36_ccff_tail;
  wire [0:19] cbx_1__1__36_chanx_left_out;
  wire [0:19] cbx_1__1__36_chanx_right_out;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__37_ccff_tail;
  wire [0:19] cbx_1__1__37_chanx_left_out;
  wire [0:19] cbx_1__1__37_chanx_right_out;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__38_ccff_tail;
  wire [0:19] cbx_1__1__38_chanx_left_out;
  wire [0:19] cbx_1__1__38_chanx_right_out;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__39_ccff_tail;
  wire [0:19] cbx_1__1__39_chanx_left_out;
  wire [0:19] cbx_1__1__39_chanx_right_out;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__3_ccff_tail;
  wire [0:19] cbx_1__1__3_chanx_left_out;
  wire [0:19] cbx_1__1__3_chanx_right_out;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__40_ccff_tail;
  wire [0:19] cbx_1__1__40_chanx_left_out;
  wire [0:19] cbx_1__1__40_chanx_right_out;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__41_ccff_tail;
  wire [0:19] cbx_1__1__41_chanx_left_out;
  wire [0:19] cbx_1__1__41_chanx_right_out;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__42_ccff_tail;
  wire [0:19] cbx_1__1__42_chanx_left_out;
  wire [0:19] cbx_1__1__42_chanx_right_out;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__43_ccff_tail;
  wire [0:19] cbx_1__1__43_chanx_left_out;
  wire [0:19] cbx_1__1__43_chanx_right_out;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__44_ccff_tail;
  wire [0:19] cbx_1__1__44_chanx_left_out;
  wire [0:19] cbx_1__1__44_chanx_right_out;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__45_ccff_tail;
  wire [0:19] cbx_1__1__45_chanx_left_out;
  wire [0:19] cbx_1__1__45_chanx_right_out;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__46_ccff_tail;
  wire [0:19] cbx_1__1__46_chanx_left_out;
  wire [0:19] cbx_1__1__46_chanx_right_out;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__47_ccff_tail;
  wire [0:19] cbx_1__1__47_chanx_left_out;
  wire [0:19] cbx_1__1__47_chanx_right_out;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__48_ccff_tail;
  wire [0:19] cbx_1__1__48_chanx_left_out;
  wire [0:19] cbx_1__1__48_chanx_right_out;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__49_ccff_tail;
  wire [0:19] cbx_1__1__49_chanx_left_out;
  wire [0:19] cbx_1__1__49_chanx_right_out;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__4_ccff_tail;
  wire [0:19] cbx_1__1__4_chanx_left_out;
  wire [0:19] cbx_1__1__4_chanx_right_out;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__50_ccff_tail;
  wire [0:19] cbx_1__1__50_chanx_left_out;
  wire [0:19] cbx_1__1__50_chanx_right_out;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__51_ccff_tail;
  wire [0:19] cbx_1__1__51_chanx_left_out;
  wire [0:19] cbx_1__1__51_chanx_right_out;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__52_ccff_tail;
  wire [0:19] cbx_1__1__52_chanx_left_out;
  wire [0:19] cbx_1__1__52_chanx_right_out;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__53_ccff_tail;
  wire [0:19] cbx_1__1__53_chanx_left_out;
  wire [0:19] cbx_1__1__53_chanx_right_out;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__54_ccff_tail;
  wire [0:19] cbx_1__1__54_chanx_left_out;
  wire [0:19] cbx_1__1__54_chanx_right_out;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__55_ccff_tail;
  wire [0:19] cbx_1__1__55_chanx_left_out;
  wire [0:19] cbx_1__1__55_chanx_right_out;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__56_ccff_tail;
  wire [0:19] cbx_1__1__56_chanx_left_out;
  wire [0:19] cbx_1__1__56_chanx_right_out;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__57_ccff_tail;
  wire [0:19] cbx_1__1__57_chanx_left_out;
  wire [0:19] cbx_1__1__57_chanx_right_out;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__58_ccff_tail;
  wire [0:19] cbx_1__1__58_chanx_left_out;
  wire [0:19] cbx_1__1__58_chanx_right_out;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__59_ccff_tail;
  wire [0:19] cbx_1__1__59_chanx_left_out;
  wire [0:19] cbx_1__1__59_chanx_right_out;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__5_ccff_tail;
  wire [0:19] cbx_1__1__5_chanx_left_out;
  wire [0:19] cbx_1__1__5_chanx_right_out;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__60_ccff_tail;
  wire [0:19] cbx_1__1__60_chanx_left_out;
  wire [0:19] cbx_1__1__60_chanx_right_out;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__61_ccff_tail;
  wire [0:19] cbx_1__1__61_chanx_left_out;
  wire [0:19] cbx_1__1__61_chanx_right_out;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__62_ccff_tail;
  wire [0:19] cbx_1__1__62_chanx_left_out;
  wire [0:19] cbx_1__1__62_chanx_right_out;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__63_ccff_tail;
  wire [0:19] cbx_1__1__63_chanx_left_out;
  wire [0:19] cbx_1__1__63_chanx_right_out;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__64_ccff_tail;
  wire [0:19] cbx_1__1__64_chanx_left_out;
  wire [0:19] cbx_1__1__64_chanx_right_out;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__65_ccff_tail;
  wire [0:19] cbx_1__1__65_chanx_left_out;
  wire [0:19] cbx_1__1__65_chanx_right_out;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__66_ccff_tail;
  wire [0:19] cbx_1__1__66_chanx_left_out;
  wire [0:19] cbx_1__1__66_chanx_right_out;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__67_ccff_tail;
  wire [0:19] cbx_1__1__67_chanx_left_out;
  wire [0:19] cbx_1__1__67_chanx_right_out;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__68_ccff_tail;
  wire [0:19] cbx_1__1__68_chanx_left_out;
  wire [0:19] cbx_1__1__68_chanx_right_out;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__69_ccff_tail;
  wire [0:19] cbx_1__1__69_chanx_left_out;
  wire [0:19] cbx_1__1__69_chanx_right_out;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__6_ccff_tail;
  wire [0:19] cbx_1__1__6_chanx_left_out;
  wire [0:19] cbx_1__1__6_chanx_right_out;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__70_ccff_tail;
  wire [0:19] cbx_1__1__70_chanx_left_out;
  wire [0:19] cbx_1__1__70_chanx_right_out;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__71_ccff_tail;
  wire [0:19] cbx_1__1__71_chanx_left_out;
  wire [0:19] cbx_1__1__71_chanx_right_out;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__72_ccff_tail;
  wire [0:19] cbx_1__1__72_chanx_left_out;
  wire [0:19] cbx_1__1__72_chanx_right_out;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__73_ccff_tail;
  wire [0:19] cbx_1__1__73_chanx_left_out;
  wire [0:19] cbx_1__1__73_chanx_right_out;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__74_ccff_tail;
  wire [0:19] cbx_1__1__74_chanx_left_out;
  wire [0:19] cbx_1__1__74_chanx_right_out;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__75_ccff_tail;
  wire [0:19] cbx_1__1__75_chanx_left_out;
  wire [0:19] cbx_1__1__75_chanx_right_out;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__76_ccff_tail;
  wire [0:19] cbx_1__1__76_chanx_left_out;
  wire [0:19] cbx_1__1__76_chanx_right_out;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__77_ccff_tail;
  wire [0:19] cbx_1__1__77_chanx_left_out;
  wire [0:19] cbx_1__1__77_chanx_right_out;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__78_ccff_tail;
  wire [0:19] cbx_1__1__78_chanx_left_out;
  wire [0:19] cbx_1__1__78_chanx_right_out;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__79_ccff_tail;
  wire [0:19] cbx_1__1__79_chanx_left_out;
  wire [0:19] cbx_1__1__79_chanx_right_out;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__7_ccff_tail;
  wire [0:19] cbx_1__1__7_chanx_left_out;
  wire [0:19] cbx_1__1__7_chanx_right_out;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__80_ccff_tail;
  wire [0:19] cbx_1__1__80_chanx_left_out;
  wire [0:19] cbx_1__1__80_chanx_right_out;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__81_ccff_tail;
  wire [0:19] cbx_1__1__81_chanx_left_out;
  wire [0:19] cbx_1__1__81_chanx_right_out;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__82_ccff_tail;
  wire [0:19] cbx_1__1__82_chanx_left_out;
  wire [0:19] cbx_1__1__82_chanx_right_out;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__83_ccff_tail;
  wire [0:19] cbx_1__1__83_chanx_left_out;
  wire [0:19] cbx_1__1__83_chanx_right_out;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__84_ccff_tail;
  wire [0:19] cbx_1__1__84_chanx_left_out;
  wire [0:19] cbx_1__1__84_chanx_right_out;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__85_ccff_tail;
  wire [0:19] cbx_1__1__85_chanx_left_out;
  wire [0:19] cbx_1__1__85_chanx_right_out;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__86_ccff_tail;
  wire [0:19] cbx_1__1__86_chanx_left_out;
  wire [0:19] cbx_1__1__86_chanx_right_out;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__87_ccff_tail;
  wire [0:19] cbx_1__1__87_chanx_left_out;
  wire [0:19] cbx_1__1__87_chanx_right_out;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__88_ccff_tail;
  wire [0:19] cbx_1__1__88_chanx_left_out;
  wire [0:19] cbx_1__1__88_chanx_right_out;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__89_ccff_tail;
  wire [0:19] cbx_1__1__89_chanx_left_out;
  wire [0:19] cbx_1__1__89_chanx_right_out;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__8_ccff_tail;
  wire [0:19] cbx_1__1__8_chanx_left_out;
  wire [0:19] cbx_1__1__8_chanx_right_out;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__90_ccff_tail;
  wire [0:19] cbx_1__1__90_chanx_left_out;
  wire [0:19] cbx_1__1__90_chanx_right_out;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__91_ccff_tail;
  wire [0:19] cbx_1__1__91_chanx_left_out;
  wire [0:19] cbx_1__1__91_chanx_right_out;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__92_ccff_tail;
  wire [0:19] cbx_1__1__92_chanx_left_out;
  wire [0:19] cbx_1__1__92_chanx_right_out;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__93_ccff_tail;
  wire [0:19] cbx_1__1__93_chanx_left_out;
  wire [0:19] cbx_1__1__93_chanx_right_out;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__94_ccff_tail;
  wire [0:19] cbx_1__1__94_chanx_left_out;
  wire [0:19] cbx_1__1__94_chanx_right_out;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__95_ccff_tail;
  wire [0:19] cbx_1__1__95_chanx_left_out;
  wire [0:19] cbx_1__1__95_chanx_right_out;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__96_ccff_tail;
  wire [0:19] cbx_1__1__96_chanx_left_out;
  wire [0:19] cbx_1__1__96_chanx_right_out;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__97_ccff_tail;
  wire [0:19] cbx_1__1__97_chanx_left_out;
  wire [0:19] cbx_1__1__97_chanx_right_out;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__98_ccff_tail;
  wire [0:19] cbx_1__1__98_chanx_left_out;
  wire [0:19] cbx_1__1__98_chanx_right_out;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__99_ccff_tail;
  wire [0:19] cbx_1__1__99_chanx_left_out;
  wire [0:19] cbx_1__1__99_chanx_right_out;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_;
  wire [0:0] cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
  wire [0:0] cbx_1__1__9_ccff_tail;
  wire [0:19] cbx_1__1__9_chanx_left_out;
  wire [0:19] cbx_1__1__9_chanx_right_out;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__0_ccff_tail;
  wire [0:19] cbx_1__3__0_chanx_left_out;
  wire [0:19] cbx_1__3__0_chanx_right_out;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__10_ccff_tail;
  wire [0:19] cbx_1__3__10_chanx_left_out;
  wire [0:19] cbx_1__3__10_chanx_right_out;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__11_ccff_tail;
  wire [0:19] cbx_1__3__11_chanx_left_out;
  wire [0:19] cbx_1__3__11_chanx_right_out;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__1_ccff_tail;
  wire [0:19] cbx_1__3__1_chanx_left_out;
  wire [0:19] cbx_1__3__1_chanx_right_out;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__2_ccff_tail;
  wire [0:19] cbx_1__3__2_chanx_left_out;
  wire [0:19] cbx_1__3__2_chanx_right_out;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__3_ccff_tail;
  wire [0:19] cbx_1__3__3_chanx_left_out;
  wire [0:19] cbx_1__3__3_chanx_right_out;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__4_ccff_tail;
  wire [0:19] cbx_1__3__4_chanx_left_out;
  wire [0:19] cbx_1__3__4_chanx_right_out;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__5_ccff_tail;
  wire [0:19] cbx_1__3__5_chanx_left_out;
  wire [0:19] cbx_1__3__5_chanx_right_out;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__6_ccff_tail;
  wire [0:19] cbx_1__3__6_chanx_left_out;
  wire [0:19] cbx_1__3__6_chanx_right_out;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__7_ccff_tail;
  wire [0:19] cbx_1__3__7_chanx_left_out;
  wire [0:19] cbx_1__3__7_chanx_right_out;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__8_ccff_tail;
  wire [0:19] cbx_1__3__8_chanx_left_out;
  wire [0:19] cbx_1__3__8_chanx_right_out;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
  wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
  wire [0:0] cbx_1__3__9_ccff_tail;
  wire [0:19] cbx_1__3__9_chanx_left_out;
  wire [0:19] cbx_1__3__9_chanx_right_out;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__0_ccff_tail;
  wire [0:19] cbx_2__3__0_chanx_left_out;
  wire [0:19] cbx_2__3__0_chanx_right_out;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__10_ccff_tail;
  wire [0:19] cbx_2__3__10_chanx_left_out;
  wire [0:19] cbx_2__3__10_chanx_right_out;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__11_ccff_tail;
  wire [0:19] cbx_2__3__11_chanx_left_out;
  wire [0:19] cbx_2__3__11_chanx_right_out;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__1_ccff_tail;
  wire [0:19] cbx_2__3__1_chanx_left_out;
  wire [0:19] cbx_2__3__1_chanx_right_out;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__2_ccff_tail;
  wire [0:19] cbx_2__3__2_chanx_left_out;
  wire [0:19] cbx_2__3__2_chanx_right_out;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__3_ccff_tail;
  wire [0:19] cbx_2__3__3_chanx_left_out;
  wire [0:19] cbx_2__3__3_chanx_right_out;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__4_ccff_tail;
  wire [0:19] cbx_2__3__4_chanx_left_out;
  wire [0:19] cbx_2__3__4_chanx_right_out;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__5_ccff_tail;
  wire [0:19] cbx_2__3__5_chanx_left_out;
  wire [0:19] cbx_2__3__5_chanx_right_out;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__6_ccff_tail;
  wire [0:19] cbx_2__3__6_chanx_left_out;
  wire [0:19] cbx_2__3__6_chanx_right_out;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__7_ccff_tail;
  wire [0:19] cbx_2__3__7_chanx_left_out;
  wire [0:19] cbx_2__3__7_chanx_right_out;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__8_ccff_tail;
  wire [0:19] cbx_2__3__8_chanx_left_out;
  wire [0:19] cbx_2__3__8_chanx_right_out;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_;
  wire [0:0] cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_;
  wire [0:0] cbx_2__3__9_ccff_tail;
  wire [0:19] cbx_2__3__9_chanx_left_out;
  wire [0:19] cbx_2__3__9_chanx_right_out;
  wire [0:0] cby_0__1__0_ccff_tail;
  wire [0:19] cby_0__1__0_chany_bottom_out;
  wire [0:19] cby_0__1__0_chany_top_out;
  wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__10_ccff_tail;
  wire [0:19] cby_0__1__10_chany_bottom_out;
  wire [0:19] cby_0__1__10_chany_top_out;
  wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__11_ccff_tail;
  wire [0:19] cby_0__1__11_chany_bottom_out;
  wire [0:19] cby_0__1__11_chany_top_out;
  wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__1_ccff_tail;
  wire [0:19] cby_0__1__1_chany_bottom_out;
  wire [0:19] cby_0__1__1_chany_top_out;
  wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__2_ccff_tail;
  wire [0:19] cby_0__1__2_chany_bottom_out;
  wire [0:19] cby_0__1__2_chany_top_out;
  wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__3_ccff_tail;
  wire [0:19] cby_0__1__3_chany_bottom_out;
  wire [0:19] cby_0__1__3_chany_top_out;
  wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__4_ccff_tail;
  wire [0:19] cby_0__1__4_chany_bottom_out;
  wire [0:19] cby_0__1__4_chany_top_out;
  wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__5_ccff_tail;
  wire [0:19] cby_0__1__5_chany_bottom_out;
  wire [0:19] cby_0__1__5_chany_top_out;
  wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__6_ccff_tail;
  wire [0:19] cby_0__1__6_chany_bottom_out;
  wire [0:19] cby_0__1__6_chany_top_out;
  wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__7_ccff_tail;
  wire [0:19] cby_0__1__7_chany_bottom_out;
  wire [0:19] cby_0__1__7_chany_top_out;
  wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__8_ccff_tail;
  wire [0:19] cby_0__1__8_chany_bottom_out;
  wire [0:19] cby_0__1__8_chany_top_out;
  wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_0__1__9_ccff_tail;
  wire [0:19] cby_0__1__9_chany_bottom_out;
  wire [0:19] cby_0__1__9_chany_top_out;
  wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__0_ccff_tail;
  wire [0:19] cby_12__1__0_chany_bottom_out;
  wire [0:19] cby_12__1__0_chany_top_out;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__1_ccff_tail;
  wire [0:19] cby_12__1__1_chany_bottom_out;
  wire [0:19] cby_12__1__1_chany_top_out;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__2_ccff_tail;
  wire [0:19] cby_12__1__2_chany_bottom_out;
  wire [0:19] cby_12__1__2_chany_top_out;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__3_ccff_tail;
  wire [0:19] cby_12__1__3_chany_bottom_out;
  wire [0:19] cby_12__1__3_chany_top_out;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__4_ccff_tail;
  wire [0:19] cby_12__1__4_chany_bottom_out;
  wire [0:19] cby_12__1__4_chany_top_out;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__5_ccff_tail;
  wire [0:19] cby_12__1__5_chany_bottom_out;
  wire [0:19] cby_12__1__5_chany_top_out;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__6_ccff_tail;
  wire [0:19] cby_12__1__6_chany_bottom_out;
  wire [0:19] cby_12__1__6_chany_top_out;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__7_ccff_tail;
  wire [0:19] cby_12__1__7_chany_bottom_out;
  wire [0:19] cby_12__1__7_chany_top_out;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__8_ccff_tail;
  wire [0:19] cby_12__1__8_chany_bottom_out;
  wire [0:19] cby_12__1__8_chany_top_out;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__1__9_ccff_tail;
  wire [0:19] cby_12__1__9_chany_bottom_out;
  wire [0:19] cby_12__1__9_chany_top_out;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_12__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__3__0_ccff_tail;
  wire [0:19] cby_12__3__0_chany_bottom_out;
  wire [0:19] cby_12__3__0_chany_top_out;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_12__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_12__3__1_ccff_tail;
  wire [0:19] cby_12__3__1_chany_bottom_out;
  wire [0:19] cby_12__3__1_chany_top_out;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_12__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
  wire [0:0] cby_1__1__0_ccff_tail;
  wire [0:19] cby_1__1__0_chany_bottom_out;
  wire [0:19] cby_1__1__0_chany_top_out;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__100_ccff_tail;
  wire [0:19] cby_1__1__100_chany_bottom_out;
  wire [0:19] cby_1__1__100_chany_top_out;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__101_ccff_tail;
  wire [0:19] cby_1__1__101_chany_bottom_out;
  wire [0:19] cby_1__1__101_chany_top_out;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__102_ccff_tail;
  wire [0:19] cby_1__1__102_chany_bottom_out;
  wire [0:19] cby_1__1__102_chany_top_out;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__103_ccff_tail;
  wire [0:19] cby_1__1__103_chany_bottom_out;
  wire [0:19] cby_1__1__103_chany_top_out;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__104_ccff_tail;
  wire [0:19] cby_1__1__104_chany_bottom_out;
  wire [0:19] cby_1__1__104_chany_top_out;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__105_ccff_tail;
  wire [0:19] cby_1__1__105_chany_bottom_out;
  wire [0:19] cby_1__1__105_chany_top_out;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__106_ccff_tail;
  wire [0:19] cby_1__1__106_chany_bottom_out;
  wire [0:19] cby_1__1__106_chany_top_out;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__107_ccff_tail;
  wire [0:19] cby_1__1__107_chany_bottom_out;
  wire [0:19] cby_1__1__107_chany_top_out;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__108_ccff_tail;
  wire [0:19] cby_1__1__108_chany_bottom_out;
  wire [0:19] cby_1__1__108_chany_top_out;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__109_ccff_tail;
  wire [0:19] cby_1__1__109_chany_bottom_out;
  wire [0:19] cby_1__1__109_chany_top_out;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__10_ccff_tail;
  wire [0:19] cby_1__1__10_chany_bottom_out;
  wire [0:19] cby_1__1__10_chany_top_out;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__11_ccff_tail;
  wire [0:19] cby_1__1__11_chany_bottom_out;
  wire [0:19] cby_1__1__11_chany_top_out;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__12_ccff_tail;
  wire [0:19] cby_1__1__12_chany_bottom_out;
  wire [0:19] cby_1__1__12_chany_top_out;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__13_ccff_tail;
  wire [0:19] cby_1__1__13_chany_bottom_out;
  wire [0:19] cby_1__1__13_chany_top_out;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__14_ccff_tail;
  wire [0:19] cby_1__1__14_chany_bottom_out;
  wire [0:19] cby_1__1__14_chany_top_out;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__15_ccff_tail;
  wire [0:19] cby_1__1__15_chany_bottom_out;
  wire [0:19] cby_1__1__15_chany_top_out;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__16_ccff_tail;
  wire [0:19] cby_1__1__16_chany_bottom_out;
  wire [0:19] cby_1__1__16_chany_top_out;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__17_ccff_tail;
  wire [0:19] cby_1__1__17_chany_bottom_out;
  wire [0:19] cby_1__1__17_chany_top_out;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__18_ccff_tail;
  wire [0:19] cby_1__1__18_chany_bottom_out;
  wire [0:19] cby_1__1__18_chany_top_out;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__19_ccff_tail;
  wire [0:19] cby_1__1__19_chany_bottom_out;
  wire [0:19] cby_1__1__19_chany_top_out;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__1_ccff_tail;
  wire [0:19] cby_1__1__1_chany_bottom_out;
  wire [0:19] cby_1__1__1_chany_top_out;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__20_ccff_tail;
  wire [0:19] cby_1__1__20_chany_bottom_out;
  wire [0:19] cby_1__1__20_chany_top_out;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__21_ccff_tail;
  wire [0:19] cby_1__1__21_chany_bottom_out;
  wire [0:19] cby_1__1__21_chany_top_out;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__22_ccff_tail;
  wire [0:19] cby_1__1__22_chany_bottom_out;
  wire [0:19] cby_1__1__22_chany_top_out;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__23_ccff_tail;
  wire [0:19] cby_1__1__23_chany_bottom_out;
  wire [0:19] cby_1__1__23_chany_top_out;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__24_ccff_tail;
  wire [0:19] cby_1__1__24_chany_bottom_out;
  wire [0:19] cby_1__1__24_chany_top_out;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__25_ccff_tail;
  wire [0:19] cby_1__1__25_chany_bottom_out;
  wire [0:19] cby_1__1__25_chany_top_out;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__26_ccff_tail;
  wire [0:19] cby_1__1__26_chany_bottom_out;
  wire [0:19] cby_1__1__26_chany_top_out;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__27_ccff_tail;
  wire [0:19] cby_1__1__27_chany_bottom_out;
  wire [0:19] cby_1__1__27_chany_top_out;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__28_ccff_tail;
  wire [0:19] cby_1__1__28_chany_bottom_out;
  wire [0:19] cby_1__1__28_chany_top_out;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__29_ccff_tail;
  wire [0:19] cby_1__1__29_chany_bottom_out;
  wire [0:19] cby_1__1__29_chany_top_out;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__2_ccff_tail;
  wire [0:19] cby_1__1__2_chany_bottom_out;
  wire [0:19] cby_1__1__2_chany_top_out;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__30_ccff_tail;
  wire [0:19] cby_1__1__30_chany_bottom_out;
  wire [0:19] cby_1__1__30_chany_top_out;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__31_ccff_tail;
  wire [0:19] cby_1__1__31_chany_bottom_out;
  wire [0:19] cby_1__1__31_chany_top_out;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__32_ccff_tail;
  wire [0:19] cby_1__1__32_chany_bottom_out;
  wire [0:19] cby_1__1__32_chany_top_out;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__33_ccff_tail;
  wire [0:19] cby_1__1__33_chany_bottom_out;
  wire [0:19] cby_1__1__33_chany_top_out;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__34_ccff_tail;
  wire [0:19] cby_1__1__34_chany_bottom_out;
  wire [0:19] cby_1__1__34_chany_top_out;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__35_ccff_tail;
  wire [0:19] cby_1__1__35_chany_bottom_out;
  wire [0:19] cby_1__1__35_chany_top_out;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__36_ccff_tail;
  wire [0:19] cby_1__1__36_chany_bottom_out;
  wire [0:19] cby_1__1__36_chany_top_out;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__37_ccff_tail;
  wire [0:19] cby_1__1__37_chany_bottom_out;
  wire [0:19] cby_1__1__37_chany_top_out;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__38_ccff_tail;
  wire [0:19] cby_1__1__38_chany_bottom_out;
  wire [0:19] cby_1__1__38_chany_top_out;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__39_ccff_tail;
  wire [0:19] cby_1__1__39_chany_bottom_out;
  wire [0:19] cby_1__1__39_chany_top_out;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__3_ccff_tail;
  wire [0:19] cby_1__1__3_chany_bottom_out;
  wire [0:19] cby_1__1__3_chany_top_out;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__40_ccff_tail;
  wire [0:19] cby_1__1__40_chany_bottom_out;
  wire [0:19] cby_1__1__40_chany_top_out;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__41_ccff_tail;
  wire [0:19] cby_1__1__41_chany_bottom_out;
  wire [0:19] cby_1__1__41_chany_top_out;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__42_ccff_tail;
  wire [0:19] cby_1__1__42_chany_bottom_out;
  wire [0:19] cby_1__1__42_chany_top_out;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__43_ccff_tail;
  wire [0:19] cby_1__1__43_chany_bottom_out;
  wire [0:19] cby_1__1__43_chany_top_out;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__44_ccff_tail;
  wire [0:19] cby_1__1__44_chany_bottom_out;
  wire [0:19] cby_1__1__44_chany_top_out;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__45_ccff_tail;
  wire [0:19] cby_1__1__45_chany_bottom_out;
  wire [0:19] cby_1__1__45_chany_top_out;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__46_ccff_tail;
  wire [0:19] cby_1__1__46_chany_bottom_out;
  wire [0:19] cby_1__1__46_chany_top_out;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__47_ccff_tail;
  wire [0:19] cby_1__1__47_chany_bottom_out;
  wire [0:19] cby_1__1__47_chany_top_out;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__48_ccff_tail;
  wire [0:19] cby_1__1__48_chany_bottom_out;
  wire [0:19] cby_1__1__48_chany_top_out;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__49_ccff_tail;
  wire [0:19] cby_1__1__49_chany_bottom_out;
  wire [0:19] cby_1__1__49_chany_top_out;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__4_ccff_tail;
  wire [0:19] cby_1__1__4_chany_bottom_out;
  wire [0:19] cby_1__1__4_chany_top_out;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__50_ccff_tail;
  wire [0:19] cby_1__1__50_chany_bottom_out;
  wire [0:19] cby_1__1__50_chany_top_out;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__51_ccff_tail;
  wire [0:19] cby_1__1__51_chany_bottom_out;
  wire [0:19] cby_1__1__51_chany_top_out;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__52_ccff_tail;
  wire [0:19] cby_1__1__52_chany_bottom_out;
  wire [0:19] cby_1__1__52_chany_top_out;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__53_ccff_tail;
  wire [0:19] cby_1__1__53_chany_bottom_out;
  wire [0:19] cby_1__1__53_chany_top_out;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__54_ccff_tail;
  wire [0:19] cby_1__1__54_chany_bottom_out;
  wire [0:19] cby_1__1__54_chany_top_out;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__55_ccff_tail;
  wire [0:19] cby_1__1__55_chany_bottom_out;
  wire [0:19] cby_1__1__55_chany_top_out;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__56_ccff_tail;
  wire [0:19] cby_1__1__56_chany_bottom_out;
  wire [0:19] cby_1__1__56_chany_top_out;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__57_ccff_tail;
  wire [0:19] cby_1__1__57_chany_bottom_out;
  wire [0:19] cby_1__1__57_chany_top_out;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__58_ccff_tail;
  wire [0:19] cby_1__1__58_chany_bottom_out;
  wire [0:19] cby_1__1__58_chany_top_out;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__59_ccff_tail;
  wire [0:19] cby_1__1__59_chany_bottom_out;
  wire [0:19] cby_1__1__59_chany_top_out;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__5_ccff_tail;
  wire [0:19] cby_1__1__5_chany_bottom_out;
  wire [0:19] cby_1__1__5_chany_top_out;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__60_ccff_tail;
  wire [0:19] cby_1__1__60_chany_bottom_out;
  wire [0:19] cby_1__1__60_chany_top_out;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__61_ccff_tail;
  wire [0:19] cby_1__1__61_chany_bottom_out;
  wire [0:19] cby_1__1__61_chany_top_out;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__62_ccff_tail;
  wire [0:19] cby_1__1__62_chany_bottom_out;
  wire [0:19] cby_1__1__62_chany_top_out;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__63_ccff_tail;
  wire [0:19] cby_1__1__63_chany_bottom_out;
  wire [0:19] cby_1__1__63_chany_top_out;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__64_ccff_tail;
  wire [0:19] cby_1__1__64_chany_bottom_out;
  wire [0:19] cby_1__1__64_chany_top_out;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__65_ccff_tail;
  wire [0:19] cby_1__1__65_chany_bottom_out;
  wire [0:19] cby_1__1__65_chany_top_out;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__66_ccff_tail;
  wire [0:19] cby_1__1__66_chany_bottom_out;
  wire [0:19] cby_1__1__66_chany_top_out;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__67_ccff_tail;
  wire [0:19] cby_1__1__67_chany_bottom_out;
  wire [0:19] cby_1__1__67_chany_top_out;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__68_ccff_tail;
  wire [0:19] cby_1__1__68_chany_bottom_out;
  wire [0:19] cby_1__1__68_chany_top_out;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__69_ccff_tail;
  wire [0:19] cby_1__1__69_chany_bottom_out;
  wire [0:19] cby_1__1__69_chany_top_out;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__6_ccff_tail;
  wire [0:19] cby_1__1__6_chany_bottom_out;
  wire [0:19] cby_1__1__6_chany_top_out;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__70_ccff_tail;
  wire [0:19] cby_1__1__70_chany_bottom_out;
  wire [0:19] cby_1__1__70_chany_top_out;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__71_ccff_tail;
  wire [0:19] cby_1__1__71_chany_bottom_out;
  wire [0:19] cby_1__1__71_chany_top_out;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__72_ccff_tail;
  wire [0:19] cby_1__1__72_chany_bottom_out;
  wire [0:19] cby_1__1__72_chany_top_out;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__73_ccff_tail;
  wire [0:19] cby_1__1__73_chany_bottom_out;
  wire [0:19] cby_1__1__73_chany_top_out;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__74_ccff_tail;
  wire [0:19] cby_1__1__74_chany_bottom_out;
  wire [0:19] cby_1__1__74_chany_top_out;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__75_ccff_tail;
  wire [0:19] cby_1__1__75_chany_bottom_out;
  wire [0:19] cby_1__1__75_chany_top_out;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__76_ccff_tail;
  wire [0:19] cby_1__1__76_chany_bottom_out;
  wire [0:19] cby_1__1__76_chany_top_out;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__77_ccff_tail;
  wire [0:19] cby_1__1__77_chany_bottom_out;
  wire [0:19] cby_1__1__77_chany_top_out;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__78_ccff_tail;
  wire [0:19] cby_1__1__78_chany_bottom_out;
  wire [0:19] cby_1__1__78_chany_top_out;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__79_ccff_tail;
  wire [0:19] cby_1__1__79_chany_bottom_out;
  wire [0:19] cby_1__1__79_chany_top_out;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__7_ccff_tail;
  wire [0:19] cby_1__1__7_chany_bottom_out;
  wire [0:19] cby_1__1__7_chany_top_out;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__80_ccff_tail;
  wire [0:19] cby_1__1__80_chany_bottom_out;
  wire [0:19] cby_1__1__80_chany_top_out;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__81_ccff_tail;
  wire [0:19] cby_1__1__81_chany_bottom_out;
  wire [0:19] cby_1__1__81_chany_top_out;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__82_ccff_tail;
  wire [0:19] cby_1__1__82_chany_bottom_out;
  wire [0:19] cby_1__1__82_chany_top_out;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__83_ccff_tail;
  wire [0:19] cby_1__1__83_chany_bottom_out;
  wire [0:19] cby_1__1__83_chany_top_out;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__84_ccff_tail;
  wire [0:19] cby_1__1__84_chany_bottom_out;
  wire [0:19] cby_1__1__84_chany_top_out;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__85_ccff_tail;
  wire [0:19] cby_1__1__85_chany_bottom_out;
  wire [0:19] cby_1__1__85_chany_top_out;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__86_ccff_tail;
  wire [0:19] cby_1__1__86_chany_bottom_out;
  wire [0:19] cby_1__1__86_chany_top_out;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__87_ccff_tail;
  wire [0:19] cby_1__1__87_chany_bottom_out;
  wire [0:19] cby_1__1__87_chany_top_out;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__88_ccff_tail;
  wire [0:19] cby_1__1__88_chany_bottom_out;
  wire [0:19] cby_1__1__88_chany_top_out;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__89_ccff_tail;
  wire [0:19] cby_1__1__89_chany_bottom_out;
  wire [0:19] cby_1__1__89_chany_top_out;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__8_ccff_tail;
  wire [0:19] cby_1__1__8_chany_bottom_out;
  wire [0:19] cby_1__1__8_chany_top_out;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__90_ccff_tail;
  wire [0:19] cby_1__1__90_chany_bottom_out;
  wire [0:19] cby_1__1__90_chany_top_out;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__91_ccff_tail;
  wire [0:19] cby_1__1__91_chany_bottom_out;
  wire [0:19] cby_1__1__91_chany_top_out;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__92_ccff_tail;
  wire [0:19] cby_1__1__92_chany_bottom_out;
  wire [0:19] cby_1__1__92_chany_top_out;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__93_ccff_tail;
  wire [0:19] cby_1__1__93_chany_bottom_out;
  wire [0:19] cby_1__1__93_chany_top_out;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__94_ccff_tail;
  wire [0:19] cby_1__1__94_chany_bottom_out;
  wire [0:19] cby_1__1__94_chany_top_out;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__95_ccff_tail;
  wire [0:19] cby_1__1__95_chany_bottom_out;
  wire [0:19] cby_1__1__95_chany_top_out;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__96_ccff_tail;
  wire [0:19] cby_1__1__96_chany_bottom_out;
  wire [0:19] cby_1__1__96_chany_top_out;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__97_ccff_tail;
  wire [0:19] cby_1__1__97_chany_bottom_out;
  wire [0:19] cby_1__1__97_chany_top_out;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__98_ccff_tail;
  wire [0:19] cby_1__1__98_chany_bottom_out;
  wire [0:19] cby_1__1__98_chany_top_out;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__99_ccff_tail;
  wire [0:19] cby_1__1__99_chany_bottom_out;
  wire [0:19] cby_1__1__99_chany_top_out;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:0] cby_1__1__9_ccff_tail;
  wire [0:19] cby_1__1__9_chany_bottom_out;
  wire [0:19] cby_1__1__9_chany_top_out;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
  wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
  wire [0:19] cby_1__3__0_chany_bottom_out;
  wire [0:19] cby_1__3__0_chany_top_out;
  wire [0:19] cby_1__3__10_chany_bottom_out;
  wire [0:19] cby_1__3__10_chany_top_out;
  wire [0:19] cby_1__3__11_chany_bottom_out;
  wire [0:19] cby_1__3__11_chany_top_out;
  wire [0:19] cby_1__3__1_chany_bottom_out;
  wire [0:19] cby_1__3__1_chany_top_out;
  wire [0:19] cby_1__3__2_chany_bottom_out;
  wire [0:19] cby_1__3__2_chany_top_out;
  wire [0:19] cby_1__3__3_chany_bottom_out;
  wire [0:19] cby_1__3__3_chany_top_out;
  wire [0:19] cby_1__3__4_chany_bottom_out;
  wire [0:19] cby_1__3__4_chany_top_out;
  wire [0:19] cby_1__3__5_chany_bottom_out;
  wire [0:19] cby_1__3__5_chany_top_out;
  wire [0:19] cby_1__3__6_chany_bottom_out;
  wire [0:19] cby_1__3__6_chany_top_out;
  wire [0:19] cby_1__3__7_chany_bottom_out;
  wire [0:19] cby_1__3__7_chany_top_out;
  wire [0:19] cby_1__3__8_chany_bottom_out;
  wire [0:19] cby_1__3__8_chany_top_out;
  wire [0:19] cby_1__3__9_chany_bottom_out;
  wire [0:19] cby_1__3__9_chany_top_out;
  wire [0:0] cby_2__3__0_ccff_tail;
  wire [0:19] cby_2__3__0_chany_bottom_out;
  wire [0:19] cby_2__3__0_chany_top_out;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__1_ccff_tail;
  wire [0:19] cby_2__3__1_chany_bottom_out;
  wire [0:19] cby_2__3__1_chany_top_out;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__2_ccff_tail;
  wire [0:19] cby_2__3__2_chany_bottom_out;
  wire [0:19] cby_2__3__2_chany_top_out;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__3_ccff_tail;
  wire [0:19] cby_2__3__3_chany_bottom_out;
  wire [0:19] cby_2__3__3_chany_top_out;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__4_ccff_tail;
  wire [0:19] cby_2__3__4_chany_bottom_out;
  wire [0:19] cby_2__3__4_chany_top_out;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__5_ccff_tail;
  wire [0:19] cby_2__3__5_chany_bottom_out;
  wire [0:19] cby_2__3__5_chany_top_out;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__6_ccff_tail;
  wire [0:19] cby_2__3__6_chany_bottom_out;
  wire [0:19] cby_2__3__6_chany_top_out;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__7_ccff_tail;
  wire [0:19] cby_2__3__7_chany_bottom_out;
  wire [0:19] cby_2__3__7_chany_top_out;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__8_ccff_tail;
  wire [0:19] cby_2__3__8_chany_bottom_out;
  wire [0:19] cby_2__3__8_chany_top_out;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] cby_2__3__9_ccff_tail;
  wire [0:19] cby_2__3__9_chany_bottom_out;
  wire [0:19] cby_2__3__9_chany_top_out;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_;
  wire [0:0] cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_;
  wire [0:0] direct_interc_0_out;
  wire [0:0] direct_interc_100_out;
  wire [0:0] direct_interc_101_out;
  wire [0:0] direct_interc_102_out;
  wire [0:0] direct_interc_103_out;
  wire [0:0] direct_interc_104_out;
  wire [0:0] direct_interc_105_out;
  wire [0:0] direct_interc_106_out;
  wire [0:0] direct_interc_107_out;
  wire [0:0] direct_interc_108_out;
  wire [0:0] direct_interc_109_out;
  wire [0:0] direct_interc_10_out;
  wire [0:0] direct_interc_110_out;
  wire [0:0] direct_interc_111_out;
  wire [0:0] direct_interc_112_out;
  wire [0:0] direct_interc_113_out;
  wire [0:0] direct_interc_114_out;
  wire [0:0] direct_interc_115_out;
  wire [0:0] direct_interc_116_out;
  wire [0:0] direct_interc_117_out;
  wire [0:0] direct_interc_118_out;
  wire [0:0] direct_interc_119_out;
  wire [0:0] direct_interc_11_out;
  wire [0:0] direct_interc_120_out;
  wire [0:0] direct_interc_121_out;
  wire [0:0] direct_interc_122_out;
  wire [0:0] direct_interc_123_out;
  wire [0:0] direct_interc_124_out;
  wire [0:0] direct_interc_125_out;
  wire [0:0] direct_interc_126_out;
  wire [0:0] direct_interc_127_out;
  wire [0:0] direct_interc_128_out;
  wire [0:0] direct_interc_129_out;
  wire [0:0] direct_interc_12_out;
  wire [0:0] direct_interc_130_out;
  wire [0:0] direct_interc_131_out;
  wire [0:0] direct_interc_132_out;
  wire [0:0] direct_interc_133_out;
  wire [0:0] direct_interc_134_out;
  wire [0:0] direct_interc_135_out;
  wire [0:0] direct_interc_136_out;
  wire [0:0] direct_interc_137_out;
  wire [0:0] direct_interc_138_out;
  wire [0:0] direct_interc_139_out;
  wire [0:0] direct_interc_13_out;
  wire [0:0] direct_interc_140_out;
  wire [0:0] direct_interc_141_out;
  wire [0:0] direct_interc_142_out;
  wire [0:0] direct_interc_143_out;
  wire [0:0] direct_interc_144_out;
  wire [0:0] direct_interc_145_out;
  wire [0:0] direct_interc_146_out;
  wire [0:0] direct_interc_147_out;
  wire [0:0] direct_interc_148_out;
  wire [0:0] direct_interc_149_out;
  wire [0:0] direct_interc_14_out;
  wire [0:0] direct_interc_150_out;
  wire [0:0] direct_interc_151_out;
  wire [0:0] direct_interc_152_out;
  wire [0:0] direct_interc_153_out;
  wire [0:0] direct_interc_154_out;
  wire [0:0] direct_interc_155_out;
  wire [0:0] direct_interc_156_out;
  wire [0:0] direct_interc_157_out;
  wire [0:0] direct_interc_158_out;
  wire [0:0] direct_interc_159_out;
  wire [0:0] direct_interc_15_out;
  wire [0:0] direct_interc_160_out;
  wire [0:0] direct_interc_161_out;
  wire [0:0] direct_interc_162_out;
  wire [0:0] direct_interc_163_out;
  wire [0:0] direct_interc_164_out;
  wire [0:0] direct_interc_165_out;
  wire [0:0] direct_interc_166_out;
  wire [0:0] direct_interc_167_out;
  wire [0:0] direct_interc_168_out;
  wire [0:0] direct_interc_169_out;
  wire [0:0] direct_interc_16_out;
  wire [0:0] direct_interc_170_out;
  wire [0:0] direct_interc_171_out;
  wire [0:0] direct_interc_172_out;
  wire [0:0] direct_interc_173_out;
  wire [0:0] direct_interc_174_out;
  wire [0:0] direct_interc_175_out;
  wire [0:0] direct_interc_176_out;
  wire [0:0] direct_interc_177_out;
  wire [0:0] direct_interc_178_out;
  wire [0:0] direct_interc_17_out;
  wire [0:0] direct_interc_18_out;
  wire [0:0] direct_interc_19_out;
  wire [0:0] direct_interc_1_out;
  wire [0:0] direct_interc_20_out;
  wire [0:0] direct_interc_21_out;
  wire [0:0] direct_interc_22_out;
  wire [0:0] direct_interc_23_out;
  wire [0:0] direct_interc_24_out;
  wire [0:0] direct_interc_25_out;
  wire [0:0] direct_interc_26_out;
  wire [0:0] direct_interc_27_out;
  wire [0:0] direct_interc_28_out;
  wire [0:0] direct_interc_29_out;
  wire [0:0] direct_interc_2_out;
  wire [0:0] direct_interc_30_out;
  wire [0:0] direct_interc_31_out;
  wire [0:0] direct_interc_32_out;
  wire [0:0] direct_interc_33_out;
  wire [0:0] direct_interc_34_out;
  wire [0:0] direct_interc_35_out;
  wire [0:0] direct_interc_36_out;
  wire [0:0] direct_interc_37_out;
  wire [0:0] direct_interc_38_out;
  wire [0:0] direct_interc_39_out;
  wire [0:0] direct_interc_3_out;
  wire [0:0] direct_interc_40_out;
  wire [0:0] direct_interc_41_out;
  wire [0:0] direct_interc_42_out;
  wire [0:0] direct_interc_43_out;
  wire [0:0] direct_interc_44_out;
  wire [0:0] direct_interc_45_out;
  wire [0:0] direct_interc_46_out;
  wire [0:0] direct_interc_47_out;
  wire [0:0] direct_interc_48_out;
  wire [0:0] direct_interc_49_out;
  wire [0:0] direct_interc_4_out;
  wire [0:0] direct_interc_50_out;
  wire [0:0] direct_interc_51_out;
  wire [0:0] direct_interc_52_out;
  wire [0:0] direct_interc_53_out;
  wire [0:0] direct_interc_54_out;
  wire [0:0] direct_interc_55_out;
  wire [0:0] direct_interc_56_out;
  wire [0:0] direct_interc_57_out;
  wire [0:0] direct_interc_58_out;
  wire [0:0] direct_interc_59_out;
  wire [0:0] direct_interc_5_out;
  wire [0:0] direct_interc_60_out;
  wire [0:0] direct_interc_61_out;
  wire [0:0] direct_interc_62_out;
  wire [0:0] direct_interc_63_out;
  wire [0:0] direct_interc_64_out;
  wire [0:0] direct_interc_65_out;
  wire [0:0] direct_interc_66_out;
  wire [0:0] direct_interc_67_out;
  wire [0:0] direct_interc_68_out;
  wire [0:0] direct_interc_69_out;
  wire [0:0] direct_interc_6_out;
  wire [0:0] direct_interc_70_out;
  wire [0:0] direct_interc_71_out;
  wire [0:0] direct_interc_72_out;
  wire [0:0] direct_interc_73_out;
  wire [0:0] direct_interc_74_out;
  wire [0:0] direct_interc_75_out;
  wire [0:0] direct_interc_76_out;
  wire [0:0] direct_interc_77_out;
  wire [0:0] direct_interc_78_out;
  wire [0:0] direct_interc_79_out;
  wire [0:0] direct_interc_7_out;
  wire [0:0] direct_interc_80_out;
  wire [0:0] direct_interc_81_out;
  wire [0:0] direct_interc_82_out;
  wire [0:0] direct_interc_83_out;
  wire [0:0] direct_interc_84_out;
  wire [0:0] direct_interc_85_out;
  wire [0:0] direct_interc_86_out;
  wire [0:0] direct_interc_87_out;
  wire [0:0] direct_interc_88_out;
  wire [0:0] direct_interc_89_out;
  wire [0:0] direct_interc_8_out;
  wire [0:0] direct_interc_90_out;
  wire [0:0] direct_interc_91_out;
  wire [0:0] direct_interc_92_out;
  wire [0:0] direct_interc_93_out;
  wire [0:0] direct_interc_94_out;
  wire [0:0] direct_interc_95_out;
  wire [0:0] direct_interc_96_out;
  wire [0:0] direct_interc_97_out;
  wire [0:0] direct_interc_98_out;
  wire [0:0] direct_interc_99_out;
  wire [0:0] direct_interc_9_out;
  wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_0_ccff_tail;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_100_ccff_tail;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_101_ccff_tail;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_102_ccff_tail;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_103_ccff_tail;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_104_ccff_tail;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_105_ccff_tail;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_106_ccff_tail;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_107_ccff_tail;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_108_ccff_tail;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_109_ccff_tail;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_10_ccff_tail;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_110_ccff_tail;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_111_ccff_tail;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_112_ccff_tail;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_113_ccff_tail;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_114_ccff_tail;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_115_ccff_tail;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_116_ccff_tail;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_117_ccff_tail;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_118_ccff_tail;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_119_ccff_tail;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_11_ccff_tail;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_12_ccff_tail;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_13_ccff_tail;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_14_ccff_tail;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_15_ccff_tail;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_16_ccff_tail;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_17_ccff_tail;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_18_ccff_tail;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_19_ccff_tail;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_1_ccff_tail;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_20_ccff_tail;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_21_ccff_tail;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_22_ccff_tail;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_23_ccff_tail;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_24_ccff_tail;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_25_ccff_tail;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_26_ccff_tail;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_27_ccff_tail;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_28_ccff_tail;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_29_ccff_tail;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_2__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_2_ccff_tail;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_30_ccff_tail;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_31_ccff_tail;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_32_ccff_tail;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_33_ccff_tail;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_34_ccff_tail;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_35_ccff_tail;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_36_ccff_tail;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_37_ccff_tail;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_38_ccff_tail;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_39_ccff_tail;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_3_ccff_tail;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_40_ccff_tail;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_41_ccff_tail;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_42_ccff_tail;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_43_ccff_tail;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_44_ccff_tail;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_45_ccff_tail;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_46_ccff_tail;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_47_ccff_tail;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_48_ccff_tail;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_49_ccff_tail;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_4_ccff_tail;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_50_ccff_tail;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_51_ccff_tail;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_52_ccff_tail;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_53_ccff_tail;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_54_ccff_tail;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_55_ccff_tail;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_56_ccff_tail;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_57_ccff_tail;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_58_ccff_tail;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_59_ccff_tail;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_5_ccff_tail;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_60_ccff_tail;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_61_ccff_tail;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_62_ccff_tail;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_63_ccff_tail;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_64_ccff_tail;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_65_ccff_tail;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_66_ccff_tail;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_67_ccff_tail;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_68_ccff_tail;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_69_ccff_tail;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_6_ccff_tail;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_70_ccff_tail;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_71_ccff_tail;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_72_ccff_tail;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_73_ccff_tail;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_74_ccff_tail;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_75_ccff_tail;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_76_ccff_tail;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_77_ccff_tail;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_78_ccff_tail;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_79_ccff_tail;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_7_ccff_tail;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_80_ccff_tail;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_81_ccff_tail;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_82_ccff_tail;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_83_ccff_tail;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_84_ccff_tail;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_85_ccff_tail;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_86_ccff_tail;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_87_ccff_tail;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_88_ccff_tail;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_89_ccff_tail;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_8__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_8_ccff_tail;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_90_ccff_tail;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_91_ccff_tail;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_92_ccff_tail;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_93_ccff_tail;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_94_ccff_tail;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_95_ccff_tail;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_96_ccff_tail;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_97_ccff_tail;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_98_ccff_tail;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_99_ccff_tail;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
  wire [0:0] grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
  wire [0:0] grid_clb_9_ccff_tail;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper;
  wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_ccff_tail;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
  wire [0:0] grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_0_ccff_tail;
  wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_10_ccff_tail;
  wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_11_ccff_tail;
  wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_1_ccff_tail;
  wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_2_ccff_tail;
  wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_3_ccff_tail;
  wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_4_ccff_tail;
  wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_5_ccff_tail;
  wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_6_ccff_tail;
  wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_7_ccff_tail;
  wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_8_ccff_tail;
  wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_left_left_9_ccff_tail;
  wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_0_ccff_tail;
  wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_10_ccff_tail;
  wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_11_ccff_tail;
  wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_1_ccff_tail;
  wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_2_ccff_tail;
  wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_3_ccff_tail;
  wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_4_ccff_tail;
  wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_5_ccff_tail;
  wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_6_ccff_tail;
  wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_7_ccff_tail;
  wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_8_ccff_tail;
  wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_right_right_9_ccff_tail;
  wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_0_ccff_tail;
  wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_10_ccff_tail;
  wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_11_ccff_tail;
  wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_1_ccff_tail;
  wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_2_ccff_tail;
  wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_3_ccff_tail;
  wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_4_ccff_tail;
  wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_5_ccff_tail;
  wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_6_ccff_tail;
  wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_7_ccff_tail;
  wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_8_ccff_tail;
  wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
  wire [0:0] grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
  wire [0:0] grid_io_top_top_9_ccff_tail;
  wire [0:0] grid_mult_18_0_ccff_tail;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_10_ccff_tail;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_11_ccff_tail;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_1_ccff_tail;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_2_ccff_tail;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_3_ccff_tail;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_4_ccff_tail;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_5_ccff_tail;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_6_ccff_tail;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_7_ccff_tail;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_8_ccff_tail;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] grid_mult_18_9_ccff_tail;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower;
  wire [0:0] grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower;
  wire [0:0] grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower;
  wire [0:0] grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper;
  wire [0:0] sb_0__0__0_ccff_tail;
  wire [0:19] sb_0__0__0_chanx_right_out;
  wire [0:19] sb_0__0__0_chany_top_out;
  wire [0:0] sb_0__12__0_ccff_tail;
  wire [0:19] sb_0__12__0_chanx_right_out;
  wire [0:19] sb_0__12__0_chany_bottom_out;
  wire [0:0] sb_0__1__0_ccff_tail;
  wire [0:19] sb_0__1__0_chanx_right_out;
  wire [0:19] sb_0__1__0_chany_bottom_out;
  wire [0:19] sb_0__1__0_chany_top_out;
  wire [0:0] sb_0__1__1_ccff_tail;
  wire [0:19] sb_0__1__1_chanx_right_out;
  wire [0:19] sb_0__1__1_chany_bottom_out;
  wire [0:19] sb_0__1__1_chany_top_out;
  wire [0:0] sb_0__1__2_ccff_tail;
  wire [0:19] sb_0__1__2_chanx_right_out;
  wire [0:19] sb_0__1__2_chany_bottom_out;
  wire [0:19] sb_0__1__2_chany_top_out;
  wire [0:0] sb_0__1__3_ccff_tail;
  wire [0:19] sb_0__1__3_chanx_right_out;
  wire [0:19] sb_0__1__3_chany_bottom_out;
  wire [0:19] sb_0__1__3_chany_top_out;
  wire [0:0] sb_0__1__4_ccff_tail;
  wire [0:19] sb_0__1__4_chanx_right_out;
  wire [0:19] sb_0__1__4_chany_bottom_out;
  wire [0:19] sb_0__1__4_chany_top_out;
  wire [0:0] sb_0__1__5_ccff_tail;
  wire [0:19] sb_0__1__5_chanx_right_out;
  wire [0:19] sb_0__1__5_chany_bottom_out;
  wire [0:19] sb_0__1__5_chany_top_out;
  wire [0:0] sb_0__1__6_ccff_tail;
  wire [0:19] sb_0__1__6_chanx_right_out;
  wire [0:19] sb_0__1__6_chany_bottom_out;
  wire [0:19] sb_0__1__6_chany_top_out;
  wire [0:0] sb_0__1__7_ccff_tail;
  wire [0:19] sb_0__1__7_chanx_right_out;
  wire [0:19] sb_0__1__7_chany_bottom_out;
  wire [0:19] sb_0__1__7_chany_top_out;
  wire [0:0] sb_0__1__8_ccff_tail;
  wire [0:19] sb_0__1__8_chanx_right_out;
  wire [0:19] sb_0__1__8_chany_bottom_out;
  wire [0:19] sb_0__1__8_chany_top_out;
  wire [0:0] sb_0__3__0_ccff_tail;
  wire [0:19] sb_0__3__0_chanx_right_out;
  wire [0:19] sb_0__3__0_chany_bottom_out;
  wire [0:19] sb_0__3__0_chany_top_out;
  wire [0:0] sb_0__3__1_ccff_tail;
  wire [0:19] sb_0__3__1_chanx_right_out;
  wire [0:19] sb_0__3__1_chany_bottom_out;
  wire [0:19] sb_0__3__1_chany_top_out;
  wire [0:19] sb_12__0__0_chanx_left_out;
  wire [0:19] sb_12__0__0_chany_top_out;
  wire [0:0] sb_12__12__0_ccff_tail;
  wire [0:19] sb_12__12__0_chanx_left_out;
  wire [0:19] sb_12__12__0_chany_bottom_out;
  wire [0:19] sb_12__1__0_chanx_left_out;
  wire [0:19] sb_12__1__0_chany_bottom_out;
  wire [0:19] sb_12__1__0_chany_top_out;
  wire [0:19] sb_12__1__1_chanx_left_out;
  wire [0:19] sb_12__1__1_chany_bottom_out;
  wire [0:19] sb_12__1__1_chany_top_out;
  wire [0:19] sb_12__1__2_chanx_left_out;
  wire [0:19] sb_12__1__2_chany_bottom_out;
  wire [0:19] sb_12__1__2_chany_top_out;
  wire [0:19] sb_12__1__3_chanx_left_out;
  wire [0:19] sb_12__1__3_chany_bottom_out;
  wire [0:19] sb_12__1__3_chany_top_out;
  wire [0:19] sb_12__1__4_chanx_left_out;
  wire [0:19] sb_12__1__4_chany_bottom_out;
  wire [0:19] sb_12__1__4_chany_top_out;
  wire [0:19] sb_12__1__5_chanx_left_out;
  wire [0:19] sb_12__1__5_chany_bottom_out;
  wire [0:19] sb_12__1__5_chany_top_out;
  wire [0:19] sb_12__1__6_chanx_left_out;
  wire [0:19] sb_12__1__6_chany_bottom_out;
  wire [0:19] sb_12__1__6_chany_top_out;
  wire [0:19] sb_12__2__0_chanx_left_out;
  wire [0:19] sb_12__2__0_chany_bottom_out;
  wire [0:19] sb_12__2__0_chany_top_out;
  wire [0:19] sb_12__2__1_chanx_left_out;
  wire [0:19] sb_12__2__1_chany_bottom_out;
  wire [0:19] sb_12__2__1_chany_top_out;
  wire [0:19] sb_12__3__0_chanx_left_out;
  wire [0:19] sb_12__3__0_chany_bottom_out;
  wire [0:19] sb_12__3__0_chany_top_out;
  wire [0:19] sb_12__3__1_chanx_left_out;
  wire [0:19] sb_12__3__1_chany_bottom_out;
  wire [0:19] sb_12__3__1_chany_top_out;
  wire [0:0] sb_1__0__0_ccff_tail;
  wire [0:19] sb_1__0__0_chanx_left_out;
  wire [0:19] sb_1__0__0_chanx_right_out;
  wire [0:19] sb_1__0__0_chany_top_out;
  wire [0:0] sb_1__0__10_ccff_tail;
  wire [0:19] sb_1__0__10_chanx_left_out;
  wire [0:19] sb_1__0__10_chanx_right_out;
  wire [0:19] sb_1__0__10_chany_top_out;
  wire [0:0] sb_1__0__1_ccff_tail;
  wire [0:19] sb_1__0__1_chanx_left_out;
  wire [0:19] sb_1__0__1_chanx_right_out;
  wire [0:19] sb_1__0__1_chany_top_out;
  wire [0:0] sb_1__0__2_ccff_tail;
  wire [0:19] sb_1__0__2_chanx_left_out;
  wire [0:19] sb_1__0__2_chanx_right_out;
  wire [0:19] sb_1__0__2_chany_top_out;
  wire [0:0] sb_1__0__3_ccff_tail;
  wire [0:19] sb_1__0__3_chanx_left_out;
  wire [0:19] sb_1__0__3_chanx_right_out;
  wire [0:19] sb_1__0__3_chany_top_out;
  wire [0:0] sb_1__0__4_ccff_tail;
  wire [0:19] sb_1__0__4_chanx_left_out;
  wire [0:19] sb_1__0__4_chanx_right_out;
  wire [0:19] sb_1__0__4_chany_top_out;
  wire [0:0] sb_1__0__5_ccff_tail;
  wire [0:19] sb_1__0__5_chanx_left_out;
  wire [0:19] sb_1__0__5_chanx_right_out;
  wire [0:19] sb_1__0__5_chany_top_out;
  wire [0:0] sb_1__0__6_ccff_tail;
  wire [0:19] sb_1__0__6_chanx_left_out;
  wire [0:19] sb_1__0__6_chanx_right_out;
  wire [0:19] sb_1__0__6_chany_top_out;
  wire [0:0] sb_1__0__7_ccff_tail;
  wire [0:19] sb_1__0__7_chanx_left_out;
  wire [0:19] sb_1__0__7_chanx_right_out;
  wire [0:19] sb_1__0__7_chany_top_out;
  wire [0:0] sb_1__0__8_ccff_tail;
  wire [0:19] sb_1__0__8_chanx_left_out;
  wire [0:19] sb_1__0__8_chanx_right_out;
  wire [0:19] sb_1__0__8_chany_top_out;
  wire [0:0] sb_1__0__9_ccff_tail;
  wire [0:19] sb_1__0__9_chanx_left_out;
  wire [0:19] sb_1__0__9_chanx_right_out;
  wire [0:19] sb_1__0__9_chany_top_out;
  wire [0:0] sb_1__12__0_ccff_tail;
  wire [0:19] sb_1__12__0_chanx_left_out;
  wire [0:19] sb_1__12__0_chanx_right_out;
  wire [0:19] sb_1__12__0_chany_bottom_out;
  wire [0:0] sb_1__12__10_ccff_tail;
  wire [0:19] sb_1__12__10_chanx_left_out;
  wire [0:19] sb_1__12__10_chanx_right_out;
  wire [0:19] sb_1__12__10_chany_bottom_out;
  wire [0:0] sb_1__12__1_ccff_tail;
  wire [0:19] sb_1__12__1_chanx_left_out;
  wire [0:19] sb_1__12__1_chanx_right_out;
  wire [0:19] sb_1__12__1_chany_bottom_out;
  wire [0:0] sb_1__12__2_ccff_tail;
  wire [0:19] sb_1__12__2_chanx_left_out;
  wire [0:19] sb_1__12__2_chanx_right_out;
  wire [0:19] sb_1__12__2_chany_bottom_out;
  wire [0:0] sb_1__12__3_ccff_tail;
  wire [0:19] sb_1__12__3_chanx_left_out;
  wire [0:19] sb_1__12__3_chanx_right_out;
  wire [0:19] sb_1__12__3_chany_bottom_out;
  wire [0:0] sb_1__12__4_ccff_tail;
  wire [0:19] sb_1__12__4_chanx_left_out;
  wire [0:19] sb_1__12__4_chanx_right_out;
  wire [0:19] sb_1__12__4_chany_bottom_out;
  wire [0:0] sb_1__12__5_ccff_tail;
  wire [0:19] sb_1__12__5_chanx_left_out;
  wire [0:19] sb_1__12__5_chanx_right_out;
  wire [0:19] sb_1__12__5_chany_bottom_out;
  wire [0:0] sb_1__12__6_ccff_tail;
  wire [0:19] sb_1__12__6_chanx_left_out;
  wire [0:19] sb_1__12__6_chanx_right_out;
  wire [0:19] sb_1__12__6_chany_bottom_out;
  wire [0:0] sb_1__12__7_ccff_tail;
  wire [0:19] sb_1__12__7_chanx_left_out;
  wire [0:19] sb_1__12__7_chanx_right_out;
  wire [0:19] sb_1__12__7_chany_bottom_out;
  wire [0:0] sb_1__12__8_ccff_tail;
  wire [0:19] sb_1__12__8_chanx_left_out;
  wire [0:19] sb_1__12__8_chanx_right_out;
  wire [0:19] sb_1__12__8_chany_bottom_out;
  wire [0:0] sb_1__12__9_ccff_tail;
  wire [0:19] sb_1__12__9_chanx_left_out;
  wire [0:19] sb_1__12__9_chanx_right_out;
  wire [0:19] sb_1__12__9_chany_bottom_out;
  wire [0:0] sb_1__1__0_ccff_tail;
  wire [0:19] sb_1__1__0_chanx_left_out;
  wire [0:19] sb_1__1__0_chanx_right_out;
  wire [0:19] sb_1__1__0_chany_bottom_out;
  wire [0:19] sb_1__1__0_chany_top_out;
  wire [0:0] sb_1__1__10_ccff_tail;
  wire [0:19] sb_1__1__10_chanx_left_out;
  wire [0:19] sb_1__1__10_chanx_right_out;
  wire [0:19] sb_1__1__10_chany_bottom_out;
  wire [0:19] sb_1__1__10_chany_top_out;
  wire [0:0] sb_1__1__11_ccff_tail;
  wire [0:19] sb_1__1__11_chanx_left_out;
  wire [0:19] sb_1__1__11_chanx_right_out;
  wire [0:19] sb_1__1__11_chany_bottom_out;
  wire [0:19] sb_1__1__11_chany_top_out;
  wire [0:0] sb_1__1__12_ccff_tail;
  wire [0:19] sb_1__1__12_chanx_left_out;
  wire [0:19] sb_1__1__12_chanx_right_out;
  wire [0:19] sb_1__1__12_chany_bottom_out;
  wire [0:19] sb_1__1__12_chany_top_out;
  wire [0:0] sb_1__1__13_ccff_tail;
  wire [0:19] sb_1__1__13_chanx_left_out;
  wire [0:19] sb_1__1__13_chanx_right_out;
  wire [0:19] sb_1__1__13_chany_bottom_out;
  wire [0:19] sb_1__1__13_chany_top_out;
  wire [0:0] sb_1__1__14_ccff_tail;
  wire [0:19] sb_1__1__14_chanx_left_out;
  wire [0:19] sb_1__1__14_chanx_right_out;
  wire [0:19] sb_1__1__14_chany_bottom_out;
  wire [0:19] sb_1__1__14_chany_top_out;
  wire [0:0] sb_1__1__15_ccff_tail;
  wire [0:19] sb_1__1__15_chanx_left_out;
  wire [0:19] sb_1__1__15_chanx_right_out;
  wire [0:19] sb_1__1__15_chany_bottom_out;
  wire [0:19] sb_1__1__15_chany_top_out;
  wire [0:0] sb_1__1__16_ccff_tail;
  wire [0:19] sb_1__1__16_chanx_left_out;
  wire [0:19] sb_1__1__16_chanx_right_out;
  wire [0:19] sb_1__1__16_chany_bottom_out;
  wire [0:19] sb_1__1__16_chany_top_out;
  wire [0:0] sb_1__1__17_ccff_tail;
  wire [0:19] sb_1__1__17_chanx_left_out;
  wire [0:19] sb_1__1__17_chanx_right_out;
  wire [0:19] sb_1__1__17_chany_bottom_out;
  wire [0:19] sb_1__1__17_chany_top_out;
  wire [0:0] sb_1__1__18_ccff_tail;
  wire [0:19] sb_1__1__18_chanx_left_out;
  wire [0:19] sb_1__1__18_chanx_right_out;
  wire [0:19] sb_1__1__18_chany_bottom_out;
  wire [0:19] sb_1__1__18_chany_top_out;
  wire [0:0] sb_1__1__19_ccff_tail;
  wire [0:19] sb_1__1__19_chanx_left_out;
  wire [0:19] sb_1__1__19_chanx_right_out;
  wire [0:19] sb_1__1__19_chany_bottom_out;
  wire [0:19] sb_1__1__19_chany_top_out;
  wire [0:0] sb_1__1__1_ccff_tail;
  wire [0:19] sb_1__1__1_chanx_left_out;
  wire [0:19] sb_1__1__1_chanx_right_out;
  wire [0:19] sb_1__1__1_chany_bottom_out;
  wire [0:19] sb_1__1__1_chany_top_out;
  wire [0:0] sb_1__1__20_ccff_tail;
  wire [0:19] sb_1__1__20_chanx_left_out;
  wire [0:19] sb_1__1__20_chanx_right_out;
  wire [0:19] sb_1__1__20_chany_bottom_out;
  wire [0:19] sb_1__1__20_chany_top_out;
  wire [0:0] sb_1__1__21_ccff_tail;
  wire [0:19] sb_1__1__21_chanx_left_out;
  wire [0:19] sb_1__1__21_chanx_right_out;
  wire [0:19] sb_1__1__21_chany_bottom_out;
  wire [0:19] sb_1__1__21_chany_top_out;
  wire [0:0] sb_1__1__22_ccff_tail;
  wire [0:19] sb_1__1__22_chanx_left_out;
  wire [0:19] sb_1__1__22_chanx_right_out;
  wire [0:19] sb_1__1__22_chany_bottom_out;
  wire [0:19] sb_1__1__22_chany_top_out;
  wire [0:0] sb_1__1__23_ccff_tail;
  wire [0:19] sb_1__1__23_chanx_left_out;
  wire [0:19] sb_1__1__23_chanx_right_out;
  wire [0:19] sb_1__1__23_chany_bottom_out;
  wire [0:19] sb_1__1__23_chany_top_out;
  wire [0:0] sb_1__1__24_ccff_tail;
  wire [0:19] sb_1__1__24_chanx_left_out;
  wire [0:19] sb_1__1__24_chanx_right_out;
  wire [0:19] sb_1__1__24_chany_bottom_out;
  wire [0:19] sb_1__1__24_chany_top_out;
  wire [0:0] sb_1__1__25_ccff_tail;
  wire [0:19] sb_1__1__25_chanx_left_out;
  wire [0:19] sb_1__1__25_chanx_right_out;
  wire [0:19] sb_1__1__25_chany_bottom_out;
  wire [0:19] sb_1__1__25_chany_top_out;
  wire [0:0] sb_1__1__26_ccff_tail;
  wire [0:19] sb_1__1__26_chanx_left_out;
  wire [0:19] sb_1__1__26_chanx_right_out;
  wire [0:19] sb_1__1__26_chany_bottom_out;
  wire [0:19] sb_1__1__26_chany_top_out;
  wire [0:0] sb_1__1__27_ccff_tail;
  wire [0:19] sb_1__1__27_chanx_left_out;
  wire [0:19] sb_1__1__27_chanx_right_out;
  wire [0:19] sb_1__1__27_chany_bottom_out;
  wire [0:19] sb_1__1__27_chany_top_out;
  wire [0:0] sb_1__1__28_ccff_tail;
  wire [0:19] sb_1__1__28_chanx_left_out;
  wire [0:19] sb_1__1__28_chanx_right_out;
  wire [0:19] sb_1__1__28_chany_bottom_out;
  wire [0:19] sb_1__1__28_chany_top_out;
  wire [0:0] sb_1__1__29_ccff_tail;
  wire [0:19] sb_1__1__29_chanx_left_out;
  wire [0:19] sb_1__1__29_chanx_right_out;
  wire [0:19] sb_1__1__29_chany_bottom_out;
  wire [0:19] sb_1__1__29_chany_top_out;
  wire [0:0] sb_1__1__2_ccff_tail;
  wire [0:19] sb_1__1__2_chanx_left_out;
  wire [0:19] sb_1__1__2_chanx_right_out;
  wire [0:19] sb_1__1__2_chany_bottom_out;
  wire [0:19] sb_1__1__2_chany_top_out;
  wire [0:0] sb_1__1__30_ccff_tail;
  wire [0:19] sb_1__1__30_chanx_left_out;
  wire [0:19] sb_1__1__30_chanx_right_out;
  wire [0:19] sb_1__1__30_chany_bottom_out;
  wire [0:19] sb_1__1__30_chany_top_out;
  wire [0:0] sb_1__1__31_ccff_tail;
  wire [0:19] sb_1__1__31_chanx_left_out;
  wire [0:19] sb_1__1__31_chanx_right_out;
  wire [0:19] sb_1__1__31_chany_bottom_out;
  wire [0:19] sb_1__1__31_chany_top_out;
  wire [0:0] sb_1__1__32_ccff_tail;
  wire [0:19] sb_1__1__32_chanx_left_out;
  wire [0:19] sb_1__1__32_chanx_right_out;
  wire [0:19] sb_1__1__32_chany_bottom_out;
  wire [0:19] sb_1__1__32_chany_top_out;
  wire [0:0] sb_1__1__33_ccff_tail;
  wire [0:19] sb_1__1__33_chanx_left_out;
  wire [0:19] sb_1__1__33_chanx_right_out;
  wire [0:19] sb_1__1__33_chany_bottom_out;
  wire [0:19] sb_1__1__33_chany_top_out;
  wire [0:0] sb_1__1__34_ccff_tail;
  wire [0:19] sb_1__1__34_chanx_left_out;
  wire [0:19] sb_1__1__34_chanx_right_out;
  wire [0:19] sb_1__1__34_chany_bottom_out;
  wire [0:19] sb_1__1__34_chany_top_out;
  wire [0:0] sb_1__1__35_ccff_tail;
  wire [0:19] sb_1__1__35_chanx_left_out;
  wire [0:19] sb_1__1__35_chanx_right_out;
  wire [0:19] sb_1__1__35_chany_bottom_out;
  wire [0:19] sb_1__1__35_chany_top_out;
  wire [0:0] sb_1__1__36_ccff_tail;
  wire [0:19] sb_1__1__36_chanx_left_out;
  wire [0:19] sb_1__1__36_chanx_right_out;
  wire [0:19] sb_1__1__36_chany_bottom_out;
  wire [0:19] sb_1__1__36_chany_top_out;
  wire [0:0] sb_1__1__37_ccff_tail;
  wire [0:19] sb_1__1__37_chanx_left_out;
  wire [0:19] sb_1__1__37_chanx_right_out;
  wire [0:19] sb_1__1__37_chany_bottom_out;
  wire [0:19] sb_1__1__37_chany_top_out;
  wire [0:0] sb_1__1__38_ccff_tail;
  wire [0:19] sb_1__1__38_chanx_left_out;
  wire [0:19] sb_1__1__38_chanx_right_out;
  wire [0:19] sb_1__1__38_chany_bottom_out;
  wire [0:19] sb_1__1__38_chany_top_out;
  wire [0:0] sb_1__1__39_ccff_tail;
  wire [0:19] sb_1__1__39_chanx_left_out;
  wire [0:19] sb_1__1__39_chanx_right_out;
  wire [0:19] sb_1__1__39_chany_bottom_out;
  wire [0:19] sb_1__1__39_chany_top_out;
  wire [0:0] sb_1__1__3_ccff_tail;
  wire [0:19] sb_1__1__3_chanx_left_out;
  wire [0:19] sb_1__1__3_chanx_right_out;
  wire [0:19] sb_1__1__3_chany_bottom_out;
  wire [0:19] sb_1__1__3_chany_top_out;
  wire [0:0] sb_1__1__40_ccff_tail;
  wire [0:19] sb_1__1__40_chanx_left_out;
  wire [0:19] sb_1__1__40_chanx_right_out;
  wire [0:19] sb_1__1__40_chany_bottom_out;
  wire [0:19] sb_1__1__40_chany_top_out;
  wire [0:0] sb_1__1__41_ccff_tail;
  wire [0:19] sb_1__1__41_chanx_left_out;
  wire [0:19] sb_1__1__41_chanx_right_out;
  wire [0:19] sb_1__1__41_chany_bottom_out;
  wire [0:19] sb_1__1__41_chany_top_out;
  wire [0:0] sb_1__1__42_ccff_tail;
  wire [0:19] sb_1__1__42_chanx_left_out;
  wire [0:19] sb_1__1__42_chanx_right_out;
  wire [0:19] sb_1__1__42_chany_bottom_out;
  wire [0:19] sb_1__1__42_chany_top_out;
  wire [0:0] sb_1__1__43_ccff_tail;
  wire [0:19] sb_1__1__43_chanx_left_out;
  wire [0:19] sb_1__1__43_chanx_right_out;
  wire [0:19] sb_1__1__43_chany_bottom_out;
  wire [0:19] sb_1__1__43_chany_top_out;
  wire [0:0] sb_1__1__44_ccff_tail;
  wire [0:19] sb_1__1__44_chanx_left_out;
  wire [0:19] sb_1__1__44_chanx_right_out;
  wire [0:19] sb_1__1__44_chany_bottom_out;
  wire [0:19] sb_1__1__44_chany_top_out;
  wire [0:0] sb_1__1__45_ccff_tail;
  wire [0:19] sb_1__1__45_chanx_left_out;
  wire [0:19] sb_1__1__45_chanx_right_out;
  wire [0:19] sb_1__1__45_chany_bottom_out;
  wire [0:19] sb_1__1__45_chany_top_out;
  wire [0:0] sb_1__1__46_ccff_tail;
  wire [0:19] sb_1__1__46_chanx_left_out;
  wire [0:19] sb_1__1__46_chanx_right_out;
  wire [0:19] sb_1__1__46_chany_bottom_out;
  wire [0:19] sb_1__1__46_chany_top_out;
  wire [0:0] sb_1__1__47_ccff_tail;
  wire [0:19] sb_1__1__47_chanx_left_out;
  wire [0:19] sb_1__1__47_chanx_right_out;
  wire [0:19] sb_1__1__47_chany_bottom_out;
  wire [0:19] sb_1__1__47_chany_top_out;
  wire [0:0] sb_1__1__48_ccff_tail;
  wire [0:19] sb_1__1__48_chanx_left_out;
  wire [0:19] sb_1__1__48_chanx_right_out;
  wire [0:19] sb_1__1__48_chany_bottom_out;
  wire [0:19] sb_1__1__48_chany_top_out;
  wire [0:0] sb_1__1__49_ccff_tail;
  wire [0:19] sb_1__1__49_chanx_left_out;
  wire [0:19] sb_1__1__49_chanx_right_out;
  wire [0:19] sb_1__1__49_chany_bottom_out;
  wire [0:19] sb_1__1__49_chany_top_out;
  wire [0:0] sb_1__1__4_ccff_tail;
  wire [0:19] sb_1__1__4_chanx_left_out;
  wire [0:19] sb_1__1__4_chanx_right_out;
  wire [0:19] sb_1__1__4_chany_bottom_out;
  wire [0:19] sb_1__1__4_chany_top_out;
  wire [0:0] sb_1__1__50_ccff_tail;
  wire [0:19] sb_1__1__50_chanx_left_out;
  wire [0:19] sb_1__1__50_chanx_right_out;
  wire [0:19] sb_1__1__50_chany_bottom_out;
  wire [0:19] sb_1__1__50_chany_top_out;
  wire [0:0] sb_1__1__51_ccff_tail;
  wire [0:19] sb_1__1__51_chanx_left_out;
  wire [0:19] sb_1__1__51_chanx_right_out;
  wire [0:19] sb_1__1__51_chany_bottom_out;
  wire [0:19] sb_1__1__51_chany_top_out;
  wire [0:0] sb_1__1__52_ccff_tail;
  wire [0:19] sb_1__1__52_chanx_left_out;
  wire [0:19] sb_1__1__52_chanx_right_out;
  wire [0:19] sb_1__1__52_chany_bottom_out;
  wire [0:19] sb_1__1__52_chany_top_out;
  wire [0:0] sb_1__1__53_ccff_tail;
  wire [0:19] sb_1__1__53_chanx_left_out;
  wire [0:19] sb_1__1__53_chanx_right_out;
  wire [0:19] sb_1__1__53_chany_bottom_out;
  wire [0:19] sb_1__1__53_chany_top_out;
  wire [0:0] sb_1__1__54_ccff_tail;
  wire [0:19] sb_1__1__54_chanx_left_out;
  wire [0:19] sb_1__1__54_chanx_right_out;
  wire [0:19] sb_1__1__54_chany_bottom_out;
  wire [0:19] sb_1__1__54_chany_top_out;
  wire [0:0] sb_1__1__55_ccff_tail;
  wire [0:19] sb_1__1__55_chanx_left_out;
  wire [0:19] sb_1__1__55_chanx_right_out;
  wire [0:19] sb_1__1__55_chany_bottom_out;
  wire [0:19] sb_1__1__55_chany_top_out;
  wire [0:0] sb_1__1__56_ccff_tail;
  wire [0:19] sb_1__1__56_chanx_left_out;
  wire [0:19] sb_1__1__56_chanx_right_out;
  wire [0:19] sb_1__1__56_chany_bottom_out;
  wire [0:19] sb_1__1__56_chany_top_out;
  wire [0:0] sb_1__1__57_ccff_tail;
  wire [0:19] sb_1__1__57_chanx_left_out;
  wire [0:19] sb_1__1__57_chanx_right_out;
  wire [0:19] sb_1__1__57_chany_bottom_out;
  wire [0:19] sb_1__1__57_chany_top_out;
  wire [0:0] sb_1__1__58_ccff_tail;
  wire [0:19] sb_1__1__58_chanx_left_out;
  wire [0:19] sb_1__1__58_chanx_right_out;
  wire [0:19] sb_1__1__58_chany_bottom_out;
  wire [0:19] sb_1__1__58_chany_top_out;
  wire [0:0] sb_1__1__59_ccff_tail;
  wire [0:19] sb_1__1__59_chanx_left_out;
  wire [0:19] sb_1__1__59_chanx_right_out;
  wire [0:19] sb_1__1__59_chany_bottom_out;
  wire [0:19] sb_1__1__59_chany_top_out;
  wire [0:0] sb_1__1__5_ccff_tail;
  wire [0:19] sb_1__1__5_chanx_left_out;
  wire [0:19] sb_1__1__5_chanx_right_out;
  wire [0:19] sb_1__1__5_chany_bottom_out;
  wire [0:19] sb_1__1__5_chany_top_out;
  wire [0:0] sb_1__1__60_ccff_tail;
  wire [0:19] sb_1__1__60_chanx_left_out;
  wire [0:19] sb_1__1__60_chanx_right_out;
  wire [0:19] sb_1__1__60_chany_bottom_out;
  wire [0:19] sb_1__1__60_chany_top_out;
  wire [0:0] sb_1__1__61_ccff_tail;
  wire [0:19] sb_1__1__61_chanx_left_out;
  wire [0:19] sb_1__1__61_chanx_right_out;
  wire [0:19] sb_1__1__61_chany_bottom_out;
  wire [0:19] sb_1__1__61_chany_top_out;
  wire [0:0] sb_1__1__62_ccff_tail;
  wire [0:19] sb_1__1__62_chanx_left_out;
  wire [0:19] sb_1__1__62_chanx_right_out;
  wire [0:19] sb_1__1__62_chany_bottom_out;
  wire [0:19] sb_1__1__62_chany_top_out;
  wire [0:0] sb_1__1__63_ccff_tail;
  wire [0:19] sb_1__1__63_chanx_left_out;
  wire [0:19] sb_1__1__63_chanx_right_out;
  wire [0:19] sb_1__1__63_chany_bottom_out;
  wire [0:19] sb_1__1__63_chany_top_out;
  wire [0:0] sb_1__1__64_ccff_tail;
  wire [0:19] sb_1__1__64_chanx_left_out;
  wire [0:19] sb_1__1__64_chanx_right_out;
  wire [0:19] sb_1__1__64_chany_bottom_out;
  wire [0:19] sb_1__1__64_chany_top_out;
  wire [0:0] sb_1__1__65_ccff_tail;
  wire [0:19] sb_1__1__65_chanx_left_out;
  wire [0:19] sb_1__1__65_chanx_right_out;
  wire [0:19] sb_1__1__65_chany_bottom_out;
  wire [0:19] sb_1__1__65_chany_top_out;
  wire [0:0] sb_1__1__66_ccff_tail;
  wire [0:19] sb_1__1__66_chanx_left_out;
  wire [0:19] sb_1__1__66_chanx_right_out;
  wire [0:19] sb_1__1__66_chany_bottom_out;
  wire [0:19] sb_1__1__66_chany_top_out;
  wire [0:0] sb_1__1__67_ccff_tail;
  wire [0:19] sb_1__1__67_chanx_left_out;
  wire [0:19] sb_1__1__67_chanx_right_out;
  wire [0:19] sb_1__1__67_chany_bottom_out;
  wire [0:19] sb_1__1__67_chany_top_out;
  wire [0:0] sb_1__1__68_ccff_tail;
  wire [0:19] sb_1__1__68_chanx_left_out;
  wire [0:19] sb_1__1__68_chanx_right_out;
  wire [0:19] sb_1__1__68_chany_bottom_out;
  wire [0:19] sb_1__1__68_chany_top_out;
  wire [0:0] sb_1__1__69_ccff_tail;
  wire [0:19] sb_1__1__69_chanx_left_out;
  wire [0:19] sb_1__1__69_chanx_right_out;
  wire [0:19] sb_1__1__69_chany_bottom_out;
  wire [0:19] sb_1__1__69_chany_top_out;
  wire [0:0] sb_1__1__6_ccff_tail;
  wire [0:19] sb_1__1__6_chanx_left_out;
  wire [0:19] sb_1__1__6_chanx_right_out;
  wire [0:19] sb_1__1__6_chany_bottom_out;
  wire [0:19] sb_1__1__6_chany_top_out;
  wire [0:0] sb_1__1__70_ccff_tail;
  wire [0:19] sb_1__1__70_chanx_left_out;
  wire [0:19] sb_1__1__70_chanx_right_out;
  wire [0:19] sb_1__1__70_chany_bottom_out;
  wire [0:19] sb_1__1__70_chany_top_out;
  wire [0:0] sb_1__1__71_ccff_tail;
  wire [0:19] sb_1__1__71_chanx_left_out;
  wire [0:19] sb_1__1__71_chanx_right_out;
  wire [0:19] sb_1__1__71_chany_bottom_out;
  wire [0:19] sb_1__1__71_chany_top_out;
  wire [0:0] sb_1__1__72_ccff_tail;
  wire [0:19] sb_1__1__72_chanx_left_out;
  wire [0:19] sb_1__1__72_chanx_right_out;
  wire [0:19] sb_1__1__72_chany_bottom_out;
  wire [0:19] sb_1__1__72_chany_top_out;
  wire [0:0] sb_1__1__73_ccff_tail;
  wire [0:19] sb_1__1__73_chanx_left_out;
  wire [0:19] sb_1__1__73_chanx_right_out;
  wire [0:19] sb_1__1__73_chany_bottom_out;
  wire [0:19] sb_1__1__73_chany_top_out;
  wire [0:0] sb_1__1__74_ccff_tail;
  wire [0:19] sb_1__1__74_chanx_left_out;
  wire [0:19] sb_1__1__74_chanx_right_out;
  wire [0:19] sb_1__1__74_chany_bottom_out;
  wire [0:19] sb_1__1__74_chany_top_out;
  wire [0:0] sb_1__1__75_ccff_tail;
  wire [0:19] sb_1__1__75_chanx_left_out;
  wire [0:19] sb_1__1__75_chanx_right_out;
  wire [0:19] sb_1__1__75_chany_bottom_out;
  wire [0:19] sb_1__1__75_chany_top_out;
  wire [0:0] sb_1__1__76_ccff_tail;
  wire [0:19] sb_1__1__76_chanx_left_out;
  wire [0:19] sb_1__1__76_chanx_right_out;
  wire [0:19] sb_1__1__76_chany_bottom_out;
  wire [0:19] sb_1__1__76_chany_top_out;
  wire [0:0] sb_1__1__7_ccff_tail;
  wire [0:19] sb_1__1__7_chanx_left_out;
  wire [0:19] sb_1__1__7_chanx_right_out;
  wire [0:19] sb_1__1__7_chany_bottom_out;
  wire [0:19] sb_1__1__7_chany_top_out;
  wire [0:0] sb_1__1__8_ccff_tail;
  wire [0:19] sb_1__1__8_chanx_left_out;
  wire [0:19] sb_1__1__8_chanx_right_out;
  wire [0:19] sb_1__1__8_chany_bottom_out;
  wire [0:19] sb_1__1__8_chany_top_out;
  wire [0:0] sb_1__1__9_ccff_tail;
  wire [0:19] sb_1__1__9_chanx_left_out;
  wire [0:19] sb_1__1__9_chanx_right_out;
  wire [0:19] sb_1__1__9_chany_bottom_out;
  wire [0:19] sb_1__1__9_chany_top_out;
  wire [0:0] sb_1__2__0_ccff_tail;
  wire [0:19] sb_1__2__0_chanx_left_out;
  wire [0:19] sb_1__2__0_chanx_right_out;
  wire [0:19] sb_1__2__0_chany_bottom_out;
  wire [0:19] sb_1__2__0_chany_top_out;
  wire [0:0] sb_1__2__10_ccff_tail;
  wire [0:19] sb_1__2__10_chanx_left_out;
  wire [0:19] sb_1__2__10_chanx_right_out;
  wire [0:19] sb_1__2__10_chany_bottom_out;
  wire [0:19] sb_1__2__10_chany_top_out;
  wire [0:0] sb_1__2__11_ccff_tail;
  wire [0:19] sb_1__2__11_chanx_left_out;
  wire [0:19] sb_1__2__11_chanx_right_out;
  wire [0:19] sb_1__2__11_chany_bottom_out;
  wire [0:19] sb_1__2__11_chany_top_out;
  wire [0:0] sb_1__2__1_ccff_tail;
  wire [0:19] sb_1__2__1_chanx_left_out;
  wire [0:19] sb_1__2__1_chanx_right_out;
  wire [0:19] sb_1__2__1_chany_bottom_out;
  wire [0:19] sb_1__2__1_chany_top_out;
  wire [0:0] sb_1__2__2_ccff_tail;
  wire [0:19] sb_1__2__2_chanx_left_out;
  wire [0:19] sb_1__2__2_chanx_right_out;
  wire [0:19] sb_1__2__2_chany_bottom_out;
  wire [0:19] sb_1__2__2_chany_top_out;
  wire [0:0] sb_1__2__3_ccff_tail;
  wire [0:19] sb_1__2__3_chanx_left_out;
  wire [0:19] sb_1__2__3_chanx_right_out;
  wire [0:19] sb_1__2__3_chany_bottom_out;
  wire [0:19] sb_1__2__3_chany_top_out;
  wire [0:0] sb_1__2__4_ccff_tail;
  wire [0:19] sb_1__2__4_chanx_left_out;
  wire [0:19] sb_1__2__4_chanx_right_out;
  wire [0:19] sb_1__2__4_chany_bottom_out;
  wire [0:19] sb_1__2__4_chany_top_out;
  wire [0:0] sb_1__2__5_ccff_tail;
  wire [0:19] sb_1__2__5_chanx_left_out;
  wire [0:19] sb_1__2__5_chanx_right_out;
  wire [0:19] sb_1__2__5_chany_bottom_out;
  wire [0:19] sb_1__2__5_chany_top_out;
  wire [0:0] sb_1__2__6_ccff_tail;
  wire [0:19] sb_1__2__6_chanx_left_out;
  wire [0:19] sb_1__2__6_chanx_right_out;
  wire [0:19] sb_1__2__6_chany_bottom_out;
  wire [0:19] sb_1__2__6_chany_top_out;
  wire [0:0] sb_1__2__7_ccff_tail;
  wire [0:19] sb_1__2__7_chanx_left_out;
  wire [0:19] sb_1__2__7_chanx_right_out;
  wire [0:19] sb_1__2__7_chany_bottom_out;
  wire [0:19] sb_1__2__7_chany_top_out;
  wire [0:0] sb_1__2__8_ccff_tail;
  wire [0:19] sb_1__2__8_chanx_left_out;
  wire [0:19] sb_1__2__8_chanx_right_out;
  wire [0:19] sb_1__2__8_chany_bottom_out;
  wire [0:19] sb_1__2__8_chany_top_out;
  wire [0:0] sb_1__2__9_ccff_tail;
  wire [0:19] sb_1__2__9_chanx_left_out;
  wire [0:19] sb_1__2__9_chanx_right_out;
  wire [0:19] sb_1__2__9_chany_bottom_out;
  wire [0:19] sb_1__2__9_chany_top_out;
  wire [0:0] sb_1__3__0_ccff_tail;
  wire [0:19] sb_1__3__0_chanx_left_out;
  wire [0:19] sb_1__3__0_chanx_right_out;
  wire [0:19] sb_1__3__0_chany_bottom_out;
  wire [0:19] sb_1__3__0_chany_top_out;
  wire [0:0] sb_1__3__10_ccff_tail;
  wire [0:19] sb_1__3__10_chanx_left_out;
  wire [0:19] sb_1__3__10_chanx_right_out;
  wire [0:19] sb_1__3__10_chany_bottom_out;
  wire [0:19] sb_1__3__10_chany_top_out;
  wire [0:0] sb_1__3__11_ccff_tail;
  wire [0:19] sb_1__3__11_chanx_left_out;
  wire [0:19] sb_1__3__11_chanx_right_out;
  wire [0:19] sb_1__3__11_chany_bottom_out;
  wire [0:19] sb_1__3__11_chany_top_out;
  wire [0:0] sb_1__3__1_ccff_tail;
  wire [0:19] sb_1__3__1_chanx_left_out;
  wire [0:19] sb_1__3__1_chanx_right_out;
  wire [0:19] sb_1__3__1_chany_bottom_out;
  wire [0:19] sb_1__3__1_chany_top_out;
  wire [0:0] sb_1__3__2_ccff_tail;
  wire [0:19] sb_1__3__2_chanx_left_out;
  wire [0:19] sb_1__3__2_chanx_right_out;
  wire [0:19] sb_1__3__2_chany_bottom_out;
  wire [0:19] sb_1__3__2_chany_top_out;
  wire [0:0] sb_1__3__3_ccff_tail;
  wire [0:19] sb_1__3__3_chanx_left_out;
  wire [0:19] sb_1__3__3_chanx_right_out;
  wire [0:19] sb_1__3__3_chany_bottom_out;
  wire [0:19] sb_1__3__3_chany_top_out;
  wire [0:0] sb_1__3__4_ccff_tail;
  wire [0:19] sb_1__3__4_chanx_left_out;
  wire [0:19] sb_1__3__4_chanx_right_out;
  wire [0:19] sb_1__3__4_chany_bottom_out;
  wire [0:19] sb_1__3__4_chany_top_out;
  wire [0:0] sb_1__3__5_ccff_tail;
  wire [0:19] sb_1__3__5_chanx_left_out;
  wire [0:19] sb_1__3__5_chanx_right_out;
  wire [0:19] sb_1__3__5_chany_bottom_out;
  wire [0:19] sb_1__3__5_chany_top_out;
  wire [0:0] sb_1__3__6_ccff_tail;
  wire [0:19] sb_1__3__6_chanx_left_out;
  wire [0:19] sb_1__3__6_chanx_right_out;
  wire [0:19] sb_1__3__6_chany_bottom_out;
  wire [0:19] sb_1__3__6_chany_top_out;
  wire [0:0] sb_1__3__7_ccff_tail;
  wire [0:19] sb_1__3__7_chanx_left_out;
  wire [0:19] sb_1__3__7_chanx_right_out;
  wire [0:19] sb_1__3__7_chany_bottom_out;
  wire [0:19] sb_1__3__7_chany_top_out;
  wire [0:0] sb_1__3__8_ccff_tail;
  wire [0:19] sb_1__3__8_chanx_left_out;
  wire [0:19] sb_1__3__8_chanx_right_out;
  wire [0:19] sb_1__3__8_chany_bottom_out;
  wire [0:19] sb_1__3__8_chany_top_out;
  wire [0:0] sb_1__3__9_ccff_tail;
  wire [0:19] sb_1__3__9_chanx_left_out;
  wire [0:19] sb_1__3__9_chanx_right_out;
  wire [0:19] sb_1__3__9_chany_bottom_out;
  wire [0:19] sb_1__3__9_chany_top_out;
  wire [0:0] sb_2__2__0_ccff_tail;
  wire [0:19] sb_2__2__0_chanx_left_out;
  wire [0:19] sb_2__2__0_chanx_right_out;
  wire [0:19] sb_2__2__0_chany_bottom_out;
  wire [0:19] sb_2__2__0_chany_top_out;
  wire [0:0] sb_2__2__1_ccff_tail;
  wire [0:19] sb_2__2__1_chanx_left_out;
  wire [0:19] sb_2__2__1_chanx_right_out;
  wire [0:19] sb_2__2__1_chany_bottom_out;
  wire [0:19] sb_2__2__1_chany_top_out;
  wire [0:0] sb_2__2__2_ccff_tail;
  wire [0:19] sb_2__2__2_chanx_left_out;
  wire [0:19] sb_2__2__2_chanx_right_out;
  wire [0:19] sb_2__2__2_chany_bottom_out;
  wire [0:19] sb_2__2__2_chany_top_out;
  wire [0:0] sb_2__2__3_ccff_tail;
  wire [0:19] sb_2__2__3_chanx_left_out;
  wire [0:19] sb_2__2__3_chanx_right_out;
  wire [0:19] sb_2__2__3_chany_bottom_out;
  wire [0:19] sb_2__2__3_chany_top_out;
  wire [0:0] sb_2__2__4_ccff_tail;
  wire [0:19] sb_2__2__4_chanx_left_out;
  wire [0:19] sb_2__2__4_chanx_right_out;
  wire [0:19] sb_2__2__4_chany_bottom_out;
  wire [0:19] sb_2__2__4_chany_top_out;
  wire [0:0] sb_2__2__5_ccff_tail;
  wire [0:19] sb_2__2__5_chanx_left_out;
  wire [0:19] sb_2__2__5_chanx_right_out;
  wire [0:19] sb_2__2__5_chany_bottom_out;
  wire [0:19] sb_2__2__5_chany_top_out;
  wire [0:0] sb_2__2__6_ccff_tail;
  wire [0:19] sb_2__2__6_chanx_left_out;
  wire [0:19] sb_2__2__6_chanx_right_out;
  wire [0:19] sb_2__2__6_chany_bottom_out;
  wire [0:19] sb_2__2__6_chany_top_out;
  wire [0:0] sb_2__2__7_ccff_tail;
  wire [0:19] sb_2__2__7_chanx_left_out;
  wire [0:19] sb_2__2__7_chanx_right_out;
  wire [0:19] sb_2__2__7_chany_bottom_out;
  wire [0:19] sb_2__2__7_chany_top_out;
  wire [0:0] sb_2__2__8_ccff_tail;
  wire [0:19] sb_2__2__8_chanx_left_out;
  wire [0:19] sb_2__2__8_chanx_right_out;
  wire [0:19] sb_2__2__8_chany_bottom_out;
  wire [0:19] sb_2__2__8_chany_top_out;
  wire [0:0] sb_2__2__9_ccff_tail;
  wire [0:19] sb_2__2__9_chanx_left_out;
  wire [0:19] sb_2__2__9_chanx_right_out;
  wire [0:19] sb_2__2__9_chany_bottom_out;
  wire [0:19] sb_2__2__9_chany_top_out;
  wire [0:0] sb_2__3__0_ccff_tail;
  wire [0:19] sb_2__3__0_chanx_left_out;
  wire [0:19] sb_2__3__0_chanx_right_out;
  wire [0:19] sb_2__3__0_chany_bottom_out;
  wire [0:19] sb_2__3__0_chany_top_out;
  wire [0:0] sb_2__3__1_ccff_tail;
  wire [0:19] sb_2__3__1_chanx_left_out;
  wire [0:19] sb_2__3__1_chanx_right_out;
  wire [0:19] sb_2__3__1_chany_bottom_out;
  wire [0:19] sb_2__3__1_chany_top_out;
  wire [0:0] sb_2__3__2_ccff_tail;
  wire [0:19] sb_2__3__2_chanx_left_out;
  wire [0:19] sb_2__3__2_chanx_right_out;
  wire [0:19] sb_2__3__2_chany_bottom_out;
  wire [0:19] sb_2__3__2_chany_top_out;
  wire [0:0] sb_2__3__3_ccff_tail;
  wire [0:19] sb_2__3__3_chanx_left_out;
  wire [0:19] sb_2__3__3_chanx_right_out;
  wire [0:19] sb_2__3__3_chany_bottom_out;
  wire [0:19] sb_2__3__3_chany_top_out;
  wire [0:0] sb_2__3__4_ccff_tail;
  wire [0:19] sb_2__3__4_chanx_left_out;
  wire [0:19] sb_2__3__4_chanx_right_out;
  wire [0:19] sb_2__3__4_chany_bottom_out;
  wire [0:19] sb_2__3__4_chany_top_out;
  wire [0:0] sb_2__3__5_ccff_tail;
  wire [0:19] sb_2__3__5_chanx_left_out;
  wire [0:19] sb_2__3__5_chanx_right_out;
  wire [0:19] sb_2__3__5_chany_bottom_out;
  wire [0:19] sb_2__3__5_chany_top_out;
  wire [0:0] sb_2__3__6_ccff_tail;
  wire [0:19] sb_2__3__6_chanx_left_out;
  wire [0:19] sb_2__3__6_chanx_right_out;
  wire [0:19] sb_2__3__6_chany_bottom_out;
  wire [0:19] sb_2__3__6_chany_top_out;
  wire [0:0] sb_2__3__7_ccff_tail;
  wire [0:19] sb_2__3__7_chanx_left_out;
  wire [0:19] sb_2__3__7_chanx_right_out;
  wire [0:19] sb_2__3__7_chany_bottom_out;
  wire [0:19] sb_2__3__7_chany_top_out;
  wire [0:0] sb_2__3__8_ccff_tail;
  wire [0:19] sb_2__3__8_chanx_left_out;
  wire [0:19] sb_2__3__8_chanx_right_out;
  wire [0:19] sb_2__3__8_chany_bottom_out;
  wire [0:19] sb_2__3__8_chany_top_out;
  wire [0:0] sb_2__3__9_ccff_tail;
  wire [0:19] sb_2__3__9_chanx_left_out;
  wire [0:19] sb_2__3__9_chanx_right_out;
  wire [0:19] sb_2__3__9_chany_bottom_out;
  wire [0:19] sb_2__3__9_chany_top_out;
  wire [1:0] UNCONN;
  wire [0:0] clk;
  wire [132:0] reg_in_feedthrough_wires;
  wire [132:0] reg_out__feedthrough_wires;
  wire [636:0] pResetWires;
  wire [287:0] Test_enWires;
  wire [287:0] resetWires;
  wire [312:0] sc_headWires;
  wire [636:0] config_enableWires;
  wire [624:0] prog_clk_0_wires;
  wire [251:0] prog_clk_1_wires;
  wire [135:0] prog_clk_2_wires;
  wire [100:0] prog_clk_3_wires;
  wire [143:0] clk_0_wires;
  wire [251:0] clk_1_wires;
  wire [135:0] clk_2_wires;
  wire [100:0] clk_3_wires;
  assign clk[0] = clk0;

  grid_clb
  grid_clb_1__1_
  (
    .clk_0_N_in(clk_1_wires[4]),
    .prog_clk_0_N_in(prog_clk_1_wires[4]),
    .prog_clk_0_W_out(prog_clk_0_wires[3]),
    .prog_clk_0_E_out(prog_clk_0_wires[1]),
    .prog_clk_0_S_out(prog_clk_0_wires[0]),
    .config_enable_N_in(config_enableWires[63]),
    .sc_head_S_out(sc_headWires[25]),
    .sc_head_N_in(sc_headWires[24]),
    .reset_E_in(resetWires[24]),
    .Test_en_E_in(Test_enWires[24]),
    .pReset_N_in(pResetWires[63]),
    .reg_in(reg_out__feedthrough_wires[0]),
    .cout(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_0_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_0_ccff_tail)
  );


  grid_clb
  grid_clb_1__2_
  (
    .clk_0_S_in(clk_1_wires[3]),
    .prog_clk_0_S_in(prog_clk_1_wires[3]),
    .prog_clk_0_W_out(prog_clk_0_wires[9]),
    .prog_clk_0_E_out(prog_clk_0_wires[7]),
    .prog_clk_0_S_out(prog_clk_0_wires[6]),
    .config_enable_N_in(config_enableWires[112]),
    .sc_head_S_out(sc_headWires[23]),
    .sc_head_N_in(sc_headWires[22]),
    .reset_E_in(resetWires[46]),
    .Test_en_E_in(Test_enWires[46]),
    .pReset_N_in(pResetWires[112]),
    .reg_in(reg_out__feedthrough_wires[1]),
    .reg_out(reg_in_feedthrough_wires[0]),
    .cout(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_1_ccff_tail)
  );


  grid_clb
  grid_clb_1__4_
  (
    .clk_0_S_in(clk_1_wires[10]),
    .prog_clk_0_S_in(prog_clk_1_wires[10]),
    .prog_clk_0_W_out(prog_clk_0_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[16]),
    .config_enable_N_in(config_enableWires[210]),
    .sc_head_S_out(sc_headWires[19]),
    .sc_head_N_in(sc_headWires[18]),
    .reset_E_in(resetWires[90]),
    .Test_en_E_in(Test_enWires[90]),
    .pReset_N_in(pResetWires[210]),
    .reg_in(reg_out__feedthrough_wires[3]),
    .reg_out(reg_in_feedthrough_wires[2]),
    .cout(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_1_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_2_ccff_tail)
  );


  grid_clb
  grid_clb_1__5_
  (
    .clk_0_N_in(clk_1_wires[18]),
    .prog_clk_0_N_in(prog_clk_1_wires[18]),
    .prog_clk_0_W_out(prog_clk_0_wires[24]),
    .prog_clk_0_E_out(prog_clk_0_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[21]),
    .config_enable_N_in(config_enableWires[259]),
    .sc_head_S_out(sc_headWires[17]),
    .sc_head_N_in(sc_headWires[16]),
    .reset_E_in(resetWires[112]),
    .Test_en_E_in(Test_enWires[112]),
    .pReset_N_in(pResetWires[259]),
    .reg_in(reg_out__feedthrough_wires[4]),
    .reg_out(reg_in_feedthrough_wires[3]),
    .cout(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_2_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_3_ccff_tail)
  );


  grid_clb
  grid_clb_1__6_
  (
    .clk_0_S_in(clk_1_wires[17]),
    .prog_clk_0_S_in(prog_clk_1_wires[17]),
    .prog_clk_0_W_out(prog_clk_0_wires[29]),
    .prog_clk_0_E_out(prog_clk_0_wires[27]),
    .prog_clk_0_S_out(prog_clk_0_wires[26]),
    .config_enable_N_in(config_enableWires[308]),
    .sc_head_S_out(sc_headWires[15]),
    .sc_head_N_in(sc_headWires[14]),
    .reset_E_in(resetWires[134]),
    .Test_en_E_in(Test_enWires[134]),
    .pReset_N_in(pResetWires[308]),
    .reg_in(reg_out__feedthrough_wires[5]),
    .reg_out(reg_in_feedthrough_wires[4]),
    .cout(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_3_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_4_ccff_tail)
  );


  grid_clb
  grid_clb_1__7_
  (
    .clk_0_N_in(clk_1_wires[25]),
    .prog_clk_0_N_in(prog_clk_1_wires[25]),
    .prog_clk_0_W_out(prog_clk_0_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[31]),
    .config_enable_N_in(config_enableWires[357]),
    .sc_head_S_out(sc_headWires[13]),
    .sc_head_N_in(sc_headWires[12]),
    .reset_E_in(resetWires[156]),
    .Test_en_E_in(Test_enWires[156]),
    .pReset_N_in(pResetWires[357]),
    .reg_in(reg_out__feedthrough_wires[6]),
    .reg_out(reg_in_feedthrough_wires[5]),
    .cout(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_4_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_5_ccff_tail)
  );


  grid_clb
  grid_clb_1__8_
  (
    .clk_0_S_in(clk_1_wires[24]),
    .prog_clk_0_S_in(prog_clk_1_wires[24]),
    .prog_clk_0_W_out(prog_clk_0_wires[39]),
    .prog_clk_0_E_out(prog_clk_0_wires[37]),
    .prog_clk_0_S_out(prog_clk_0_wires[36]),
    .config_enable_N_in(config_enableWires[406]),
    .sc_head_S_out(sc_headWires[11]),
    .sc_head_N_in(sc_headWires[10]),
    .reset_E_in(resetWires[178]),
    .Test_en_E_in(Test_enWires[178]),
    .pReset_N_in(pResetWires[406]),
    .reg_in(reg_out__feedthrough_wires[7]),
    .reg_out(reg_in_feedthrough_wires[6]),
    .cout(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_5_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_6_ccff_tail)
  );


  grid_clb
  grid_clb_1__9_
  (
    .clk_0_N_in(clk_1_wires[32]),
    .prog_clk_0_N_in(prog_clk_1_wires[32]),
    .prog_clk_0_W_out(prog_clk_0_wires[44]),
    .prog_clk_0_E_out(prog_clk_0_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[41]),
    .config_enable_N_in(config_enableWires[455]),
    .sc_head_S_out(sc_headWires[9]),
    .sc_head_N_in(sc_headWires[8]),
    .reset_E_in(resetWires[200]),
    .Test_en_E_in(Test_enWires[200]),
    .pReset_N_in(pResetWires[455]),
    .reg_in(reg_out__feedthrough_wires[8]),
    .reg_out(reg_in_feedthrough_wires[7]),
    .cout(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_1__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_7_ccff_tail)
  );


  grid_clb
  grid_clb_1__11_
  (
    .clk_0_N_in(clk_1_wires[39]),
    .prog_clk_0_N_in(prog_clk_1_wires[39]),
    .prog_clk_0_W_out(prog_clk_0_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[51]),
    .config_enable_N_in(config_enableWires[553]),
    .sc_head_S_out(sc_headWires[5]),
    .sc_head_N_in(sc_headWires[4]),
    .reset_E_in(resetWires[244]),
    .Test_en_E_in(Test_enWires[244]),
    .pReset_N_in(pResetWires[553]),
    .reg_in(reg_out__feedthrough_wires[10]),
    .reg_out(reg_in_feedthrough_wires[9]),
    .cout(grid_clb_1__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_6_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_8_ccff_tail)
  );


  grid_clb
  grid_clb_1__12_
  (
    .clk_0_S_in(clk_1_wires[38]),
    .prog_clk_0_S_in(prog_clk_1_wires[38]),
    .prog_clk_0_W_out(prog_clk_0_wires[61]),
    .prog_clk_0_N_out(prog_clk_0_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[56]),
    .config_enable_N_in(config_enableWires[602]),
    .sc_head_S_out(sc_headWires[3]),
    .sc_head_N_in(sc_headWires[2]),
    .reset_E_in(resetWires[266]),
    .Test_en_E_in(Test_enWires[266]),
    .pReset_N_in(pResetWires[602]),
    .reg_out(reg_in_feedthrough_wires[10]),
    .cout(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_1__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_9_ccff_tail)
  );


  grid_clb
  grid_clb_2__1_
  (
    .clk_0_N_in(clk_1_wires[6]),
    .prog_clk_0_N_in(prog_clk_1_wires[6]),
    .prog_clk_0_E_out(prog_clk_0_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[63]),
    .config_enable_N_in(config_enableWires[68]),
    .sc_head_N_out(sc_headWires[29]),
    .sc_head_S_in(sc_headWires[28]),
    .reset_W_out(resetWires[26]),
    .reset_E_in(resetWires[25]),
    .Test_en_W_out(Test_enWires[26]),
    .Test_en_E_in(Test_enWires[25]),
    .pReset_N_in(pResetWires[68]),
    .reg_in(reg_out__feedthrough_wires[11]),
    .cout(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_7_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__10_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_10_ccff_tail)
  );


  grid_clb
  grid_clb_2__2_
  (
    .clk_0_S_in(clk_1_wires[5]),
    .prog_clk_0_S_in(prog_clk_1_wires[5]),
    .prog_clk_0_E_out(prog_clk_0_wires[67]),
    .prog_clk_0_S_out(prog_clk_0_wires[66]),
    .config_enable_N_in(config_enableWires[117]),
    .sc_head_N_out(sc_headWires[31]),
    .sc_head_S_in(sc_headWires[30]),
    .reset_W_out(resetWires[48]),
    .reset_E_in(resetWires[47]),
    .Test_en_W_out(Test_enWires[48]),
    .Test_en_E_in(Test_enWires[47]),
    .pReset_N_in(pResetWires[117]),
    .reg_in(reg_out__feedthrough_wires[12]),
    .reg_out(reg_in_feedthrough_wires[11]),
    .cout(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__11_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_11_ccff_tail)
  );


  grid_clb
  grid_clb_2__4_
  (
    .clk_0_S_in(clk_1_wires[12]),
    .prog_clk_0_S_in(prog_clk_1_wires[12]),
    .prog_clk_0_E_out(prog_clk_0_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[72]),
    .config_enable_N_in(config_enableWires[215]),
    .sc_head_N_out(sc_headWires[35]),
    .sc_head_S_in(sc_headWires[34]),
    .reset_W_out(resetWires[92]),
    .reset_E_in(resetWires[91]),
    .Test_en_W_out(Test_enWires[92]),
    .Test_en_E_in(Test_enWires[91]),
    .pReset_N_in(pResetWires[215]),
    .reg_in(reg_out__feedthrough_wires[14]),
    .reg_out(reg_in_feedthrough_wires[13]),
    .cout(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_8_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__12_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_12_ccff_tail)
  );


  grid_clb
  grid_clb_2__5_
  (
    .clk_0_N_in(clk_1_wires[20]),
    .prog_clk_0_N_in(prog_clk_1_wires[20]),
    .prog_clk_0_E_out(prog_clk_0_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[75]),
    .config_enable_N_in(config_enableWires[264]),
    .sc_head_N_out(sc_headWires[37]),
    .sc_head_S_in(sc_headWires[36]),
    .reset_W_out(resetWires[114]),
    .reset_E_in(resetWires[113]),
    .Test_en_W_out(Test_enWires[114]),
    .Test_en_E_in(Test_enWires[113]),
    .pReset_N_in(pResetWires[264]),
    .reg_in(reg_out__feedthrough_wires[15]),
    .reg_out(reg_in_feedthrough_wires[14]),
    .cout(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_9_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__13_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_13_ccff_tail)
  );


  grid_clb
  grid_clb_2__6_
  (
    .clk_0_S_in(clk_1_wires[19]),
    .prog_clk_0_S_in(prog_clk_1_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[79]),
    .prog_clk_0_S_out(prog_clk_0_wires[78]),
    .config_enable_N_in(config_enableWires[313]),
    .sc_head_N_out(sc_headWires[39]),
    .sc_head_S_in(sc_headWires[38]),
    .reset_W_out(resetWires[136]),
    .reset_E_in(resetWires[135]),
    .Test_en_W_out(Test_enWires[136]),
    .Test_en_E_in(Test_enWires[135]),
    .pReset_N_in(pResetWires[313]),
    .reg_in(reg_out__feedthrough_wires[16]),
    .reg_out(reg_in_feedthrough_wires[15]),
    .cout(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_10_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__14_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_14_ccff_tail)
  );


  grid_clb
  grid_clb_2__7_
  (
    .clk_0_N_in(clk_1_wires[27]),
    .prog_clk_0_N_in(prog_clk_1_wires[27]),
    .prog_clk_0_E_out(prog_clk_0_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[81]),
    .config_enable_N_in(config_enableWires[362]),
    .sc_head_N_out(sc_headWires[41]),
    .sc_head_S_in(sc_headWires[40]),
    .reset_W_out(resetWires[158]),
    .reset_E_in(resetWires[157]),
    .Test_en_W_out(Test_enWires[158]),
    .Test_en_E_in(Test_enWires[157]),
    .pReset_N_in(pResetWires[362]),
    .reg_in(reg_out__feedthrough_wires[17]),
    .reg_out(reg_in_feedthrough_wires[16]),
    .cout(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_11_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__15_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_15_ccff_tail)
  );


  grid_clb
  grid_clb_2__8_
  (
    .clk_0_S_in(clk_1_wires[26]),
    .prog_clk_0_S_in(prog_clk_1_wires[26]),
    .prog_clk_0_E_out(prog_clk_0_wires[85]),
    .prog_clk_0_S_out(prog_clk_0_wires[84]),
    .config_enable_N_in(config_enableWires[411]),
    .sc_head_N_out(sc_headWires[43]),
    .sc_head_S_in(sc_headWires[42]),
    .reset_W_out(resetWires[180]),
    .reset_E_in(resetWires[179]),
    .Test_en_W_out(Test_enWires[180]),
    .Test_en_E_in(Test_enWires[179]),
    .pReset_N_in(pResetWires[411]),
    .reg_in(reg_out__feedthrough_wires[18]),
    .reg_out(reg_in_feedthrough_wires[17]),
    .cout(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_12_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__16_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_16_ccff_tail)
  );


  grid_clb
  grid_clb_2__9_
  (
    .clk_0_N_in(clk_1_wires[34]),
    .prog_clk_0_N_in(prog_clk_1_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[87]),
    .config_enable_N_in(config_enableWires[460]),
    .sc_head_N_out(sc_headWires[45]),
    .sc_head_S_in(sc_headWires[44]),
    .reset_W_out(resetWires[202]),
    .reset_E_in(resetWires[201]),
    .Test_en_W_out(Test_enWires[202]),
    .Test_en_E_in(Test_enWires[201]),
    .pReset_N_in(pResetWires[460]),
    .reg_in(reg_out__feedthrough_wires[19]),
    .reg_out(reg_in_feedthrough_wires[18]),
    .cout(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_2__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__17_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_17_ccff_tail)
  );


  grid_clb
  grid_clb_2__11_
  (
    .clk_0_N_in(clk_1_wires[41]),
    .prog_clk_0_N_in(prog_clk_1_wires[41]),
    .prog_clk_0_E_out(prog_clk_0_wires[94]),
    .prog_clk_0_S_out(prog_clk_0_wires[93]),
    .config_enable_N_in(config_enableWires[558]),
    .sc_head_N_out(sc_headWires[49]),
    .sc_head_S_in(sc_headWires[48]),
    .reset_W_out(resetWires[246]),
    .reset_E_in(resetWires[245]),
    .Test_en_W_out(Test_enWires[246]),
    .Test_en_E_in(Test_enWires[245]),
    .pReset_N_in(pResetWires[558]),
    .reg_in(reg_out__feedthrough_wires[21]),
    .reg_out(reg_in_feedthrough_wires[20]),
    .cout(grid_clb_2__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_13_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__18_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_18_ccff_tail)
  );


  grid_clb
  grid_clb_2__12_
  (
    .clk_0_S_in(clk_1_wires[40]),
    .prog_clk_0_S_in(prog_clk_1_wires[40]),
    .prog_clk_0_N_out(prog_clk_0_wires[99]),
    .prog_clk_0_E_out(prog_clk_0_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[96]),
    .config_enable_N_in(config_enableWires[606]),
    .sc_head_N_out(sc_headWires[51]),
    .sc_head_S_in(sc_headWires[50]),
    .reset_W_out(resetWires[268]),
    .reset_E_in(resetWires[267]),
    .Test_en_W_out(Test_enWires[268]),
    .Test_en_E_in(Test_enWires[267]),
    .pReset_N_in(pResetWires[606]),
    .reg_out(reg_in_feedthrough_wires[21]),
    .cout(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_2__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__19_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_19_ccff_tail)
  );


  grid_clb
  grid_clb_3__1_
  (
    .clk_0_N_in(clk_1_wires[46]),
    .prog_clk_0_N_in(prog_clk_1_wires[46]),
    .prog_clk_0_E_out(prog_clk_0_wires[102]),
    .prog_clk_0_S_out(prog_clk_0_wires[101]),
    .config_enable_N_in(config_enableWires[72]),
    .sc_head_S_out(sc_headWires[77]),
    .sc_head_N_in(sc_headWires[76]),
    .reset_W_out(resetWires[28]),
    .reset_E_in(resetWires[27]),
    .Test_en_W_out(Test_enWires[28]),
    .Test_en_E_in(Test_enWires[27]),
    .pReset_N_in(pResetWires[72]),
    .reg_in(reg_out__feedthrough_wires[22]),
    .cout(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_14_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__20_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_20_ccff_tail)
  );


  grid_clb
  grid_clb_3__2_
  (
    .clk_0_S_in(clk_1_wires[45]),
    .prog_clk_0_S_in(prog_clk_1_wires[45]),
    .prog_clk_0_E_out(prog_clk_0_wires[105]),
    .prog_clk_0_S_out(prog_clk_0_wires[104]),
    .config_enable_N_in(config_enableWires[121]),
    .sc_head_S_out(sc_headWires[75]),
    .sc_head_N_in(sc_headWires[74]),
    .reset_W_out(resetWires[50]),
    .reset_E_in(resetWires[49]),
    .Test_en_W_out(Test_enWires[50]),
    .Test_en_E_in(Test_enWires[49]),
    .pReset_N_in(pResetWires[121]),
    .reg_in(reg_out__feedthrough_wires[23]),
    .reg_out(reg_in_feedthrough_wires[22]),
    .cout(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__21_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_21_ccff_tail)
  );


  grid_clb
  grid_clb_3__4_
  (
    .clk_0_S_in(clk_1_wires[52]),
    .prog_clk_0_S_in(prog_clk_1_wires[52]),
    .prog_clk_0_E_out(prog_clk_0_wires[111]),
    .prog_clk_0_S_out(prog_clk_0_wires[110]),
    .config_enable_N_in(config_enableWires[219]),
    .sc_head_S_out(sc_headWires[71]),
    .sc_head_N_in(sc_headWires[70]),
    .reset_W_out(resetWires[94]),
    .reset_E_in(resetWires[93]),
    .Test_en_W_out(Test_enWires[94]),
    .Test_en_E_in(Test_enWires[93]),
    .pReset_N_in(pResetWires[219]),
    .reg_in(reg_out__feedthrough_wires[25]),
    .reg_out(reg_in_feedthrough_wires[24]),
    .cout(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_15_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__22_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_22_ccff_tail)
  );


  grid_clb
  grid_clb_3__5_
  (
    .clk_0_N_in(clk_1_wires[60]),
    .prog_clk_0_N_in(prog_clk_1_wires[60]),
    .prog_clk_0_E_out(prog_clk_0_wires[114]),
    .prog_clk_0_S_out(prog_clk_0_wires[113]),
    .config_enable_N_in(config_enableWires[268]),
    .sc_head_S_out(sc_headWires[69]),
    .sc_head_N_in(sc_headWires[68]),
    .reset_W_out(resetWires[116]),
    .reset_E_in(resetWires[115]),
    .Test_en_W_out(Test_enWires[116]),
    .Test_en_E_in(Test_enWires[115]),
    .pReset_N_in(pResetWires[268]),
    .reg_in(reg_out__feedthrough_wires[26]),
    .reg_out(reg_in_feedthrough_wires[25]),
    .cout(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_16_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__23_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_23_ccff_tail)
  );


  grid_clb
  grid_clb_3__6_
  (
    .clk_0_S_in(clk_1_wires[59]),
    .prog_clk_0_S_in(prog_clk_1_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[117]),
    .prog_clk_0_S_out(prog_clk_0_wires[116]),
    .config_enable_N_in(config_enableWires[317]),
    .sc_head_S_out(sc_headWires[67]),
    .sc_head_N_in(sc_headWires[66]),
    .reset_W_out(resetWires[138]),
    .reset_E_in(resetWires[137]),
    .Test_en_W_out(Test_enWires[138]),
    .Test_en_E_in(Test_enWires[137]),
    .pReset_N_in(pResetWires[317]),
    .reg_in(reg_out__feedthrough_wires[27]),
    .reg_out(reg_in_feedthrough_wires[26]),
    .cout(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_17_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__24_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_24_ccff_tail)
  );


  grid_clb
  grid_clb_3__7_
  (
    .clk_0_N_in(clk_1_wires[67]),
    .prog_clk_0_N_in(prog_clk_1_wires[67]),
    .prog_clk_0_E_out(prog_clk_0_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[119]),
    .config_enable_N_in(config_enableWires[366]),
    .sc_head_S_out(sc_headWires[65]),
    .sc_head_N_in(sc_headWires[64]),
    .reset_W_out(resetWires[160]),
    .reset_E_in(resetWires[159]),
    .Test_en_W_out(Test_enWires[160]),
    .Test_en_E_in(Test_enWires[159]),
    .pReset_N_in(pResetWires[366]),
    .reg_in(reg_out__feedthrough_wires[28]),
    .reg_out(reg_in_feedthrough_wires[27]),
    .cout(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_18_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__25_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_25_ccff_tail)
  );


  grid_clb
  grid_clb_3__8_
  (
    .clk_0_S_in(clk_1_wires[66]),
    .prog_clk_0_S_in(prog_clk_1_wires[66]),
    .prog_clk_0_E_out(prog_clk_0_wires[123]),
    .prog_clk_0_S_out(prog_clk_0_wires[122]),
    .config_enable_N_in(config_enableWires[415]),
    .sc_head_S_out(sc_headWires[63]),
    .sc_head_N_in(sc_headWires[62]),
    .reset_W_out(resetWires[182]),
    .reset_E_in(resetWires[181]),
    .Test_en_W_out(Test_enWires[182]),
    .Test_en_E_in(Test_enWires[181]),
    .pReset_N_in(pResetWires[415]),
    .reg_in(reg_out__feedthrough_wires[29]),
    .reg_out(reg_in_feedthrough_wires[28]),
    .cout(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_19_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__26_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_26_ccff_tail)
  );


  grid_clb
  grid_clb_3__9_
  (
    .clk_0_N_in(clk_1_wires[74]),
    .prog_clk_0_N_in(prog_clk_1_wires[74]),
    .prog_clk_0_E_out(prog_clk_0_wires[126]),
    .prog_clk_0_S_out(prog_clk_0_wires[125]),
    .config_enable_N_in(config_enableWires[464]),
    .sc_head_S_out(sc_headWires[61]),
    .sc_head_N_in(sc_headWires[60]),
    .reset_W_out(resetWires[204]),
    .reset_E_in(resetWires[203]),
    .Test_en_W_out(Test_enWires[204]),
    .Test_en_E_in(Test_enWires[203]),
    .pReset_N_in(pResetWires[464]),
    .reg_in(reg_out__feedthrough_wires[30]),
    .reg_out(reg_in_feedthrough_wires[29]),
    .cout(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_3__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__27_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_27_ccff_tail)
  );


  grid_clb
  grid_clb_3__11_
  (
    .clk_0_N_in(clk_1_wires[81]),
    .prog_clk_0_N_in(prog_clk_1_wires[81]),
    .prog_clk_0_E_out(prog_clk_0_wires[132]),
    .prog_clk_0_S_out(prog_clk_0_wires[131]),
    .config_enable_N_in(config_enableWires[562]),
    .sc_head_S_out(sc_headWires[57]),
    .sc_head_N_in(sc_headWires[56]),
    .reset_W_out(resetWires[248]),
    .reset_E_in(resetWires[247]),
    .Test_en_W_out(Test_enWires[248]),
    .Test_en_E_in(Test_enWires[247]),
    .pReset_N_in(pResetWires[562]),
    .reg_in(reg_out__feedthrough_wires[32]),
    .reg_out(reg_in_feedthrough_wires[31]),
    .cout(grid_clb_3__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_20_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__28_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_28_ccff_tail)
  );


  grid_clb
  grid_clb_3__12_
  (
    .clk_0_S_in(clk_1_wires[80]),
    .prog_clk_0_S_in(prog_clk_1_wires[80]),
    .prog_clk_0_N_out(prog_clk_0_wires[137]),
    .prog_clk_0_E_out(prog_clk_0_wires[135]),
    .prog_clk_0_S_out(prog_clk_0_wires[134]),
    .config_enable_N_in(config_enableWires[609]),
    .sc_head_S_out(sc_headWires[55]),
    .sc_head_N_in(sc_headWires[54]),
    .reset_W_out(resetWires[270]),
    .reset_E_in(resetWires[269]),
    .Test_en_W_out(Test_enWires[270]),
    .Test_en_E_in(Test_enWires[269]),
    .pReset_N_in(pResetWires[609]),
    .reg_out(reg_in_feedthrough_wires[32]),
    .cout(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_3__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__29_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_29_ccff_tail)
  );


  grid_clb
  grid_clb_4__1_
  (
    .clk_0_N_in(clk_1_wires[48]),
    .prog_clk_0_N_in(prog_clk_1_wires[48]),
    .prog_clk_0_E_out(prog_clk_0_wires[140]),
    .prog_clk_0_S_out(prog_clk_0_wires[139]),
    .config_enable_N_in(config_enableWires[76]),
    .sc_head_N_out(sc_headWires[81]),
    .sc_head_S_in(sc_headWires[80]),
    .reset_W_out(resetWires[30]),
    .reset_E_in(resetWires[29]),
    .Test_en_W_out(Test_enWires[30]),
    .Test_en_E_in(Test_enWires[29]),
    .pReset_N_in(pResetWires[76]),
    .reg_in(reg_out__feedthrough_wires[33]),
    .cout(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_21_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__30_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_30_ccff_tail)
  );


  grid_clb
  grid_clb_4__2_
  (
    .clk_0_S_in(clk_1_wires[47]),
    .prog_clk_0_S_in(prog_clk_1_wires[47]),
    .prog_clk_0_E_out(prog_clk_0_wires[143]),
    .prog_clk_0_S_out(prog_clk_0_wires[142]),
    .config_enable_N_in(config_enableWires[125]),
    .sc_head_N_out(sc_headWires[83]),
    .sc_head_S_in(sc_headWires[82]),
    .reset_W_out(resetWires[52]),
    .reset_E_in(resetWires[51]),
    .Test_en_W_out(Test_enWires[52]),
    .Test_en_E_in(Test_enWires[51]),
    .pReset_N_in(pResetWires[125]),
    .reg_in(reg_out__feedthrough_wires[34]),
    .reg_out(reg_in_feedthrough_wires[33]),
    .cout(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__31_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_31_ccff_tail)
  );


  grid_clb
  grid_clb_4__4_
  (
    .clk_0_S_in(clk_1_wires[54]),
    .prog_clk_0_S_in(prog_clk_1_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[149]),
    .prog_clk_0_S_out(prog_clk_0_wires[148]),
    .config_enable_N_in(config_enableWires[223]),
    .sc_head_N_out(sc_headWires[87]),
    .sc_head_S_in(sc_headWires[86]),
    .reset_W_out(resetWires[96]),
    .reset_E_in(resetWires[95]),
    .Test_en_W_out(Test_enWires[96]),
    .Test_en_E_in(Test_enWires[95]),
    .pReset_N_in(pResetWires[223]),
    .reg_in(reg_out__feedthrough_wires[36]),
    .reg_out(reg_in_feedthrough_wires[35]),
    .cout(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_22_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__32_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_32_ccff_tail)
  );


  grid_clb
  grid_clb_4__5_
  (
    .clk_0_N_in(clk_1_wires[62]),
    .prog_clk_0_N_in(prog_clk_1_wires[62]),
    .prog_clk_0_E_out(prog_clk_0_wires[152]),
    .prog_clk_0_S_out(prog_clk_0_wires[151]),
    .config_enable_N_in(config_enableWires[272]),
    .sc_head_N_out(sc_headWires[89]),
    .sc_head_S_in(sc_headWires[88]),
    .reset_W_out(resetWires[118]),
    .reset_E_in(resetWires[117]),
    .Test_en_W_out(Test_enWires[118]),
    .Test_en_E_in(Test_enWires[117]),
    .pReset_N_in(pResetWires[272]),
    .reg_in(reg_out__feedthrough_wires[37]),
    .reg_out(reg_in_feedthrough_wires[36]),
    .cout(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_23_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__33_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_33_ccff_tail)
  );


  grid_clb
  grid_clb_4__6_
  (
    .clk_0_S_in(clk_1_wires[61]),
    .prog_clk_0_S_in(prog_clk_1_wires[61]),
    .prog_clk_0_E_out(prog_clk_0_wires[155]),
    .prog_clk_0_S_out(prog_clk_0_wires[154]),
    .config_enable_N_in(config_enableWires[321]),
    .sc_head_N_out(sc_headWires[91]),
    .sc_head_S_in(sc_headWires[90]),
    .reset_W_out(resetWires[140]),
    .reset_E_in(resetWires[139]),
    .Test_en_W_out(Test_enWires[140]),
    .Test_en_E_in(Test_enWires[139]),
    .pReset_N_in(pResetWires[321]),
    .reg_in(reg_out__feedthrough_wires[38]),
    .reg_out(reg_in_feedthrough_wires[37]),
    .cout(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_24_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__34_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_34_ccff_tail)
  );


  grid_clb
  grid_clb_4__7_
  (
    .clk_0_N_in(clk_1_wires[69]),
    .prog_clk_0_N_in(prog_clk_1_wires[69]),
    .prog_clk_0_E_out(prog_clk_0_wires[158]),
    .prog_clk_0_S_out(prog_clk_0_wires[157]),
    .config_enable_N_in(config_enableWires[370]),
    .sc_head_N_out(sc_headWires[93]),
    .sc_head_S_in(sc_headWires[92]),
    .reset_W_out(resetWires[162]),
    .reset_E_in(resetWires[161]),
    .Test_en_W_out(Test_enWires[162]),
    .Test_en_E_in(Test_enWires[161]),
    .pReset_N_in(pResetWires[370]),
    .reg_in(reg_out__feedthrough_wires[39]),
    .reg_out(reg_in_feedthrough_wires[38]),
    .cout(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_25_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__35_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_35_ccff_tail)
  );


  grid_clb
  grid_clb_4__8_
  (
    .clk_0_S_in(clk_1_wires[68]),
    .prog_clk_0_S_in(prog_clk_1_wires[68]),
    .prog_clk_0_E_out(prog_clk_0_wires[161]),
    .prog_clk_0_S_out(prog_clk_0_wires[160]),
    .config_enable_N_in(config_enableWires[419]),
    .sc_head_N_out(sc_headWires[95]),
    .sc_head_S_in(sc_headWires[94]),
    .reset_W_out(resetWires[184]),
    .reset_E_in(resetWires[183]),
    .Test_en_W_out(Test_enWires[184]),
    .Test_en_E_in(Test_enWires[183]),
    .pReset_N_in(pResetWires[419]),
    .reg_in(reg_out__feedthrough_wires[40]),
    .reg_out(reg_in_feedthrough_wires[39]),
    .cout(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_26_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__36_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_36_ccff_tail)
  );


  grid_clb
  grid_clb_4__9_
  (
    .clk_0_N_in(clk_1_wires[76]),
    .prog_clk_0_N_in(prog_clk_1_wires[76]),
    .prog_clk_0_E_out(prog_clk_0_wires[164]),
    .prog_clk_0_S_out(prog_clk_0_wires[163]),
    .config_enable_N_in(config_enableWires[468]),
    .sc_head_N_out(sc_headWires[97]),
    .sc_head_S_in(sc_headWires[96]),
    .reset_W_out(resetWires[206]),
    .reset_E_in(resetWires[205]),
    .Test_en_W_out(Test_enWires[206]),
    .Test_en_E_in(Test_enWires[205]),
    .pReset_N_in(pResetWires[468]),
    .reg_in(reg_out__feedthrough_wires[41]),
    .reg_out(reg_in_feedthrough_wires[40]),
    .cout(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_4__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__37_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_37_ccff_tail)
  );


  grid_clb
  grid_clb_4__11_
  (
    .clk_0_N_in(clk_1_wires[83]),
    .prog_clk_0_N_in(prog_clk_1_wires[83]),
    .prog_clk_0_E_out(prog_clk_0_wires[170]),
    .prog_clk_0_S_out(prog_clk_0_wires[169]),
    .config_enable_N_in(config_enableWires[566]),
    .sc_head_N_out(sc_headWires[101]),
    .sc_head_S_in(sc_headWires[100]),
    .reset_W_out(resetWires[250]),
    .reset_E_in(resetWires[249]),
    .Test_en_W_out(Test_enWires[250]),
    .Test_en_E_in(Test_enWires[249]),
    .pReset_N_in(pResetWires[566]),
    .reg_in(reg_out__feedthrough_wires[43]),
    .reg_out(reg_in_feedthrough_wires[42]),
    .cout(grid_clb_4__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_27_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__38_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_38_ccff_tail)
  );


  grid_clb
  grid_clb_4__12_
  (
    .clk_0_S_in(clk_1_wires[82]),
    .prog_clk_0_S_in(prog_clk_1_wires[82]),
    .prog_clk_0_N_out(prog_clk_0_wires[175]),
    .prog_clk_0_E_out(prog_clk_0_wires[173]),
    .prog_clk_0_S_out(prog_clk_0_wires[172]),
    .config_enable_N_in(config_enableWires[612]),
    .sc_head_N_out(sc_headWires[103]),
    .sc_head_S_in(sc_headWires[102]),
    .reset_W_out(resetWires[272]),
    .reset_E_in(resetWires[271]),
    .Test_en_W_out(Test_enWires[272]),
    .Test_en_E_in(Test_enWires[271]),
    .pReset_N_in(pResetWires[612]),
    .reg_out(reg_in_feedthrough_wires[43]),
    .cout(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_4__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__39_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_39_ccff_tail)
  );


  grid_clb
  grid_clb_5__1_
  (
    .clk_0_N_in(clk_1_wires[88]),
    .prog_clk_0_N_in(prog_clk_1_wires[88]),
    .prog_clk_0_E_out(prog_clk_0_wires[178]),
    .prog_clk_0_S_out(prog_clk_0_wires[177]),
    .config_enable_N_in(config_enableWires[80]),
    .sc_head_S_out(sc_headWires[129]),
    .sc_head_N_in(sc_headWires[128]),
    .reset_W_out(resetWires[32]),
    .reset_E_in(resetWires[31]),
    .Test_en_W_out(Test_enWires[32]),
    .Test_en_E_in(Test_enWires[31]),
    .pReset_N_in(pResetWires[80]),
    .reg_in(reg_out__feedthrough_wires[44]),
    .cout(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_28_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__40_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_40_ccff_tail)
  );


  grid_clb
  grid_clb_5__2_
  (
    .clk_0_S_in(clk_1_wires[87]),
    .prog_clk_0_S_in(prog_clk_1_wires[87]),
    .prog_clk_0_E_out(prog_clk_0_wires[181]),
    .prog_clk_0_S_out(prog_clk_0_wires[180]),
    .config_enable_N_in(config_enableWires[129]),
    .sc_head_S_out(sc_headWires[127]),
    .sc_head_N_in(sc_headWires[126]),
    .reset_W_out(resetWires[54]),
    .reset_E_in(resetWires[53]),
    .Test_en_W_out(Test_enWires[54]),
    .Test_en_E_in(Test_enWires[53]),
    .pReset_N_in(pResetWires[129]),
    .reg_in(reg_out__feedthrough_wires[45]),
    .reg_out(reg_in_feedthrough_wires[44]),
    .cout(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__41_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_41_ccff_tail)
  );


  grid_clb
  grid_clb_5__4_
  (
    .clk_0_S_in(clk_1_wires[94]),
    .prog_clk_0_S_in(prog_clk_1_wires[94]),
    .prog_clk_0_E_out(prog_clk_0_wires[187]),
    .prog_clk_0_S_out(prog_clk_0_wires[186]),
    .config_enable_N_in(config_enableWires[227]),
    .sc_head_S_out(sc_headWires[123]),
    .sc_head_N_in(sc_headWires[122]),
    .reset_W_out(resetWires[98]),
    .reset_E_in(resetWires[97]),
    .Test_en_W_out(Test_enWires[98]),
    .Test_en_E_in(Test_enWires[97]),
    .pReset_N_in(pResetWires[227]),
    .reg_in(reg_out__feedthrough_wires[47]),
    .reg_out(reg_in_feedthrough_wires[46]),
    .cout(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_29_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__42_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_42_ccff_tail)
  );


  grid_clb
  grid_clb_5__5_
  (
    .clk_0_N_in(clk_1_wires[102]),
    .prog_clk_0_N_in(prog_clk_1_wires[102]),
    .prog_clk_0_E_out(prog_clk_0_wires[190]),
    .prog_clk_0_S_out(prog_clk_0_wires[189]),
    .config_enable_N_in(config_enableWires[276]),
    .sc_head_S_out(sc_headWires[121]),
    .sc_head_N_in(sc_headWires[120]),
    .reset_W_out(resetWires[120]),
    .reset_E_in(resetWires[119]),
    .Test_en_W_out(Test_enWires[120]),
    .Test_en_E_in(Test_enWires[119]),
    .pReset_N_in(pResetWires[276]),
    .reg_in(reg_out__feedthrough_wires[48]),
    .reg_out(reg_in_feedthrough_wires[47]),
    .cout(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_30_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__43_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_43_ccff_tail)
  );


  grid_clb
  grid_clb_5__6_
  (
    .clk_0_S_in(clk_1_wires[101]),
    .prog_clk_0_S_in(prog_clk_1_wires[101]),
    .prog_clk_0_E_out(prog_clk_0_wires[193]),
    .prog_clk_0_S_out(prog_clk_0_wires[192]),
    .config_enable_N_in(config_enableWires[325]),
    .sc_head_S_out(sc_headWires[119]),
    .sc_head_N_in(sc_headWires[118]),
    .reset_W_out(resetWires[142]),
    .reset_E_in(resetWires[141]),
    .Test_en_W_out(Test_enWires[142]),
    .Test_en_E_in(Test_enWires[141]),
    .pReset_N_in(pResetWires[325]),
    .reg_in(reg_out__feedthrough_wires[49]),
    .reg_out(reg_in_feedthrough_wires[48]),
    .cout(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_31_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__44_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_44_ccff_tail)
  );


  grid_clb
  grid_clb_5__7_
  (
    .clk_0_N_in(clk_1_wires[109]),
    .prog_clk_0_N_in(prog_clk_1_wires[109]),
    .prog_clk_0_E_out(prog_clk_0_wires[196]),
    .prog_clk_0_S_out(prog_clk_0_wires[195]),
    .config_enable_N_in(config_enableWires[374]),
    .sc_head_S_out(sc_headWires[117]),
    .sc_head_N_in(sc_headWires[116]),
    .reset_W_out(resetWires[164]),
    .reset_E_in(resetWires[163]),
    .Test_en_W_out(Test_enWires[164]),
    .Test_en_E_in(Test_enWires[163]),
    .pReset_N_in(pResetWires[374]),
    .reg_in(reg_out__feedthrough_wires[50]),
    .reg_out(reg_in_feedthrough_wires[49]),
    .cout(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_32_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__45_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_45_ccff_tail)
  );


  grid_clb
  grid_clb_5__8_
  (
    .clk_0_S_in(clk_1_wires[108]),
    .prog_clk_0_S_in(prog_clk_1_wires[108]),
    .prog_clk_0_E_out(prog_clk_0_wires[199]),
    .prog_clk_0_S_out(prog_clk_0_wires[198]),
    .config_enable_N_in(config_enableWires[423]),
    .sc_head_S_out(sc_headWires[115]),
    .sc_head_N_in(sc_headWires[114]),
    .reset_W_out(resetWires[186]),
    .reset_E_in(resetWires[185]),
    .Test_en_W_out(Test_enWires[186]),
    .Test_en_E_in(Test_enWires[185]),
    .pReset_N_in(pResetWires[423]),
    .reg_in(reg_out__feedthrough_wires[51]),
    .reg_out(reg_in_feedthrough_wires[50]),
    .cout(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_33_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__46_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_46_ccff_tail)
  );


  grid_clb
  grid_clb_5__9_
  (
    .clk_0_N_in(clk_1_wires[116]),
    .prog_clk_0_N_in(prog_clk_1_wires[116]),
    .prog_clk_0_E_out(prog_clk_0_wires[202]),
    .prog_clk_0_S_out(prog_clk_0_wires[201]),
    .config_enable_N_in(config_enableWires[472]),
    .sc_head_S_out(sc_headWires[113]),
    .sc_head_N_in(sc_headWires[112]),
    .reset_W_out(resetWires[208]),
    .reset_E_in(resetWires[207]),
    .Test_en_W_out(Test_enWires[208]),
    .Test_en_E_in(Test_enWires[207]),
    .pReset_N_in(pResetWires[472]),
    .reg_in(reg_out__feedthrough_wires[52]),
    .reg_out(reg_in_feedthrough_wires[51]),
    .cout(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_5__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__47_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_47_ccff_tail)
  );


  grid_clb
  grid_clb_5__11_
  (
    .clk_0_N_in(clk_1_wires[123]),
    .prog_clk_0_N_in(prog_clk_1_wires[123]),
    .prog_clk_0_E_out(prog_clk_0_wires[208]),
    .prog_clk_0_S_out(prog_clk_0_wires[207]),
    .config_enable_N_in(config_enableWires[570]),
    .sc_head_S_out(sc_headWires[109]),
    .sc_head_N_in(sc_headWires[108]),
    .reset_W_out(resetWires[252]),
    .reset_E_in(resetWires[251]),
    .Test_en_W_out(Test_enWires[252]),
    .Test_en_E_in(Test_enWires[251]),
    .pReset_N_in(pResetWires[570]),
    .reg_in(reg_out__feedthrough_wires[54]),
    .reg_out(reg_in_feedthrough_wires[53]),
    .cout(grid_clb_5__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_34_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__48_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_48_ccff_tail)
  );


  grid_clb
  grid_clb_5__12_
  (
    .clk_0_S_in(clk_1_wires[122]),
    .prog_clk_0_S_in(prog_clk_1_wires[122]),
    .prog_clk_0_N_out(prog_clk_0_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[211]),
    .prog_clk_0_S_out(prog_clk_0_wires[210]),
    .config_enable_N_in(config_enableWires[615]),
    .sc_head_S_out(sc_headWires[107]),
    .sc_head_N_in(sc_headWires[106]),
    .reset_W_out(resetWires[274]),
    .reset_E_in(resetWires[273]),
    .Test_en_W_out(Test_enWires[274]),
    .Test_en_E_in(Test_enWires[273]),
    .pReset_N_in(pResetWires[615]),
    .reg_out(reg_in_feedthrough_wires[54]),
    .cout(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_5__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__49_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_49_ccff_tail)
  );


  grid_clb
  grid_clb_6__1_
  (
    .clk_0_N_in(clk_1_wires[90]),
    .prog_clk_0_N_in(prog_clk_1_wires[90]),
    .prog_clk_0_E_out(prog_clk_0_wires[216]),
    .prog_clk_0_S_out(prog_clk_0_wires[215]),
    .config_enable_N_in(config_enableWires[84]),
    .sc_head_N_out(sc_headWires[133]),
    .sc_head_S_in(sc_headWires[132]),
    .reset_W_out(resetWires[34]),
    .reset_E_in(resetWires[33]),
    .Test_en_W_out(Test_enWires[34]),
    .Test_en_E_in(Test_enWires[33]),
    .pReset_N_in(pResetWires[84]),
    .reg_in(reg_out__feedthrough_wires[55]),
    .cout(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_35_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__50_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_50_ccff_tail)
  );


  grid_clb
  grid_clb_6__2_
  (
    .clk_0_S_in(clk_1_wires[89]),
    .prog_clk_0_S_in(prog_clk_1_wires[89]),
    .prog_clk_0_E_out(prog_clk_0_wires[219]),
    .prog_clk_0_S_out(prog_clk_0_wires[218]),
    .config_enable_N_in(config_enableWires[133]),
    .sc_head_N_out(sc_headWires[135]),
    .sc_head_S_in(sc_headWires[134]),
    .reset_W_out(resetWires[56]),
    .reset_E_in(resetWires[55]),
    .Test_en_W_out(Test_enWires[56]),
    .Test_en_E_in(Test_enWires[55]),
    .pReset_N_in(pResetWires[133]),
    .reg_in(reg_out__feedthrough_wires[56]),
    .reg_out(reg_in_feedthrough_wires[55]),
    .cout(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__51_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_51_ccff_tail)
  );


  grid_clb
  grid_clb_6__4_
  (
    .clk_0_S_in(clk_1_wires[96]),
    .prog_clk_0_S_in(prog_clk_1_wires[96]),
    .prog_clk_0_E_out(prog_clk_0_wires[225]),
    .prog_clk_0_S_out(prog_clk_0_wires[224]),
    .config_enable_N_in(config_enableWires[231]),
    .sc_head_N_out(sc_headWires[139]),
    .sc_head_S_in(sc_headWires[138]),
    .reset_W_out(resetWires[100]),
    .reset_E_in(resetWires[99]),
    .Test_en_W_out(Test_enWires[100]),
    .Test_en_E_in(Test_enWires[99]),
    .pReset_N_in(pResetWires[231]),
    .reg_in(reg_out__feedthrough_wires[58]),
    .reg_out(reg_in_feedthrough_wires[57]),
    .cout(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_36_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__52_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_52_ccff_tail)
  );


  grid_clb
  grid_clb_6__5_
  (
    .clk_0_N_in(clk_1_wires[104]),
    .prog_clk_0_N_in(prog_clk_1_wires[104]),
    .prog_clk_0_E_out(prog_clk_0_wires[228]),
    .prog_clk_0_S_out(prog_clk_0_wires[227]),
    .config_enable_N_in(config_enableWires[280]),
    .sc_head_N_out(sc_headWires[141]),
    .sc_head_S_in(sc_headWires[140]),
    .reset_W_out(resetWires[122]),
    .reset_E_in(resetWires[121]),
    .Test_en_W_out(Test_enWires[122]),
    .Test_en_E_in(Test_enWires[121]),
    .pReset_N_in(pResetWires[280]),
    .reg_in(reg_out__feedthrough_wires[59]),
    .reg_out(reg_in_feedthrough_wires[58]),
    .cout(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_37_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__53_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_53_ccff_tail)
  );


  grid_clb
  grid_clb_6__6_
  (
    .clk_0_S_in(clk_1_wires[103]),
    .prog_clk_0_S_in(prog_clk_1_wires[103]),
    .prog_clk_0_E_out(prog_clk_0_wires[231]),
    .prog_clk_0_S_out(prog_clk_0_wires[230]),
    .config_enable_N_in(config_enableWires[329]),
    .sc_head_N_out(sc_headWires[143]),
    .sc_head_S_in(sc_headWires[142]),
    .reset_W_out(resetWires[144]),
    .reset_E_in(resetWires[143]),
    .Test_en_W_out(Test_enWires[144]),
    .Test_en_E_in(Test_enWires[143]),
    .pReset_N_in(pResetWires[329]),
    .reg_in(reg_out__feedthrough_wires[60]),
    .reg_out(reg_in_feedthrough_wires[59]),
    .cout(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_38_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__54_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_54_ccff_tail)
  );


  grid_clb
  grid_clb_6__7_
  (
    .clk_0_N_in(clk_1_wires[111]),
    .prog_clk_0_N_in(prog_clk_1_wires[111]),
    .prog_clk_0_E_out(prog_clk_0_wires[234]),
    .prog_clk_0_S_out(prog_clk_0_wires[233]),
    .config_enable_N_in(config_enableWires[378]),
    .sc_head_N_out(sc_headWires[145]),
    .sc_head_S_in(sc_headWires[144]),
    .reset_W_out(resetWires[166]),
    .reset_E_in(resetWires[165]),
    .Test_en_W_out(Test_enWires[166]),
    .Test_en_E_in(Test_enWires[165]),
    .pReset_N_in(pResetWires[378]),
    .reg_in(reg_out__feedthrough_wires[61]),
    .reg_out(reg_in_feedthrough_wires[60]),
    .cout(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_39_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__55_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_55_ccff_tail)
  );


  grid_clb
  grid_clb_6__8_
  (
    .clk_0_S_in(clk_1_wires[110]),
    .prog_clk_0_S_in(prog_clk_1_wires[110]),
    .prog_clk_0_E_out(prog_clk_0_wires[237]),
    .prog_clk_0_S_out(prog_clk_0_wires[236]),
    .config_enable_N_in(config_enableWires[427]),
    .sc_head_N_out(sc_headWires[147]),
    .sc_head_S_in(sc_headWires[146]),
    .reset_W_out(resetWires[188]),
    .reset_E_in(resetWires[187]),
    .Test_en_W_out(Test_enWires[188]),
    .Test_en_E_in(Test_enWires[187]),
    .pReset_N_in(pResetWires[427]),
    .reg_in(reg_out__feedthrough_wires[62]),
    .reg_out(reg_in_feedthrough_wires[61]),
    .cout(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_40_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__56_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_56_ccff_tail)
  );


  grid_clb
  grid_clb_6__9_
  (
    .clk_0_N_in(clk_1_wires[118]),
    .prog_clk_0_N_in(prog_clk_1_wires[118]),
    .prog_clk_0_E_out(prog_clk_0_wires[240]),
    .prog_clk_0_S_out(prog_clk_0_wires[239]),
    .config_enable_N_in(config_enableWires[476]),
    .sc_head_N_out(sc_headWires[149]),
    .sc_head_S_in(sc_headWires[148]),
    .reset_W_out(resetWires[210]),
    .reset_E_in(resetWires[209]),
    .Test_en_W_out(Test_enWires[210]),
    .Test_en_E_in(Test_enWires[209]),
    .pReset_N_in(pResetWires[476]),
    .reg_in(reg_out__feedthrough_wires[63]),
    .reg_out(reg_in_feedthrough_wires[62]),
    .cout(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_6__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__57_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_57_ccff_tail)
  );


  grid_clb
  grid_clb_6__11_
  (
    .clk_0_N_in(clk_1_wires[125]),
    .prog_clk_0_N_in(prog_clk_1_wires[125]),
    .prog_clk_0_E_out(prog_clk_0_wires[246]),
    .prog_clk_0_S_out(prog_clk_0_wires[245]),
    .config_enable_N_in(config_enableWires[574]),
    .sc_head_N_out(sc_headWires[153]),
    .sc_head_S_in(sc_headWires[152]),
    .reset_W_out(resetWires[254]),
    .reset_E_in(resetWires[253]),
    .Test_en_W_out(Test_enWires[254]),
    .Test_en_E_in(Test_enWires[253]),
    .pReset_N_in(pResetWires[574]),
    .reg_in(reg_out__feedthrough_wires[65]),
    .reg_out(reg_in_feedthrough_wires[64]),
    .cout(grid_clb_6__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_41_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__58_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_58_ccff_tail)
  );


  grid_clb
  grid_clb_6__12_
  (
    .clk_0_S_in(clk_1_wires[124]),
    .prog_clk_0_S_in(prog_clk_1_wires[124]),
    .prog_clk_0_N_out(prog_clk_0_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[249]),
    .prog_clk_0_S_out(prog_clk_0_wires[248]),
    .config_enable_N_in(config_enableWires[618]),
    .sc_head_N_out(sc_headWires[155]),
    .sc_head_S_in(sc_headWires[154]),
    .reset_W_out(resetWires[276]),
    .reset_E_in(resetWires[275]),
    .Test_en_W_out(Test_enWires[276]),
    .Test_en_E_in(Test_enWires[275]),
    .pReset_N_in(pResetWires[618]),
    .reg_out(reg_in_feedthrough_wires[65]),
    .cout(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_6__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__59_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_59_ccff_tail)
  );


  grid_clb
  grid_clb_7__1_
  (
    .clk_0_N_in(clk_1_wires[130]),
    .prog_clk_0_N_in(prog_clk_1_wires[130]),
    .prog_clk_0_E_out(prog_clk_0_wires[254]),
    .prog_clk_0_S_out(prog_clk_0_wires[253]),
    .config_enable_N_in(config_enableWires[88]),
    .sc_head_S_out(sc_headWires[181]),
    .sc_head_N_in(sc_headWires[180]),
    .reset_E_out(resetWires[36]),
    .reset_W_in(resetWires[35]),
    .Test_en_E_out(Test_enWires[36]),
    .Test_en_W_in(Test_enWires[35]),
    .pReset_N_in(pResetWires[88]),
    .reg_in(reg_out__feedthrough_wires[66]),
    .cout(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_42_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__60_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_60_ccff_tail)
  );


  grid_clb
  grid_clb_7__2_
  (
    .clk_0_S_in(clk_1_wires[129]),
    .prog_clk_0_S_in(prog_clk_1_wires[129]),
    .prog_clk_0_E_out(prog_clk_0_wires[257]),
    .prog_clk_0_S_out(prog_clk_0_wires[256]),
    .config_enable_N_in(config_enableWires[137]),
    .sc_head_S_out(sc_headWires[179]),
    .sc_head_N_in(sc_headWires[178]),
    .reset_E_out(resetWires[58]),
    .reset_W_in(resetWires[57]),
    .Test_en_E_out(Test_enWires[58]),
    .Test_en_W_in(Test_enWires[57]),
    .pReset_N_in(pResetWires[137]),
    .reg_in(reg_out__feedthrough_wires[67]),
    .reg_out(reg_in_feedthrough_wires[66]),
    .cout(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_7__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__61_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_61_ccff_tail)
  );


  grid_clb
  grid_clb_7__4_
  (
    .clk_0_S_in(clk_1_wires[136]),
    .prog_clk_0_S_in(prog_clk_1_wires[136]),
    .prog_clk_0_E_out(prog_clk_0_wires[263]),
    .prog_clk_0_S_out(prog_clk_0_wires[262]),
    .config_enable_N_in(config_enableWires[235]),
    .sc_head_S_out(sc_headWires[175]),
    .sc_head_N_in(sc_headWires[174]),
    .reset_E_out(resetWires[102]),
    .reset_W_in(resetWires[101]),
    .Test_en_E_out(Test_enWires[102]),
    .Test_en_W_in(Test_enWires[101]),
    .pReset_N_in(pResetWires[235]),
    .reg_in(reg_out__feedthrough_wires[69]),
    .reg_out(reg_in_feedthrough_wires[68]),
    .cout(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_43_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__62_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_62_ccff_tail)
  );


  grid_clb
  grid_clb_7__5_
  (
    .clk_0_N_in(clk_1_wires[144]),
    .prog_clk_0_N_in(prog_clk_1_wires[144]),
    .prog_clk_0_E_out(prog_clk_0_wires[266]),
    .prog_clk_0_S_out(prog_clk_0_wires[265]),
    .config_enable_N_in(config_enableWires[284]),
    .sc_head_S_out(sc_headWires[173]),
    .sc_head_N_in(sc_headWires[172]),
    .reset_E_out(resetWires[124]),
    .reset_W_in(resetWires[123]),
    .Test_en_E_out(Test_enWires[124]),
    .Test_en_W_in(Test_enWires[123]),
    .pReset_N_in(pResetWires[284]),
    .reg_in(reg_out__feedthrough_wires[70]),
    .reg_out(reg_in_feedthrough_wires[69]),
    .cout(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_44_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__63_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_63_ccff_tail)
  );


  grid_clb
  grid_clb_7__6_
  (
    .clk_0_S_in(clk_1_wires[143]),
    .prog_clk_0_S_in(prog_clk_1_wires[143]),
    .prog_clk_0_E_out(prog_clk_0_wires[269]),
    .prog_clk_0_S_out(prog_clk_0_wires[268]),
    .config_enable_N_in(config_enableWires[333]),
    .sc_head_S_out(sc_headWires[171]),
    .sc_head_N_in(sc_headWires[170]),
    .reset_E_out(resetWires[146]),
    .reset_W_in(resetWires[145]),
    .Test_en_E_out(Test_enWires[146]),
    .Test_en_W_in(Test_enWires[145]),
    .pReset_N_in(pResetWires[333]),
    .reg_in(reg_out__feedthrough_wires[71]),
    .reg_out(reg_in_feedthrough_wires[70]),
    .cout(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_45_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__64_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_64_ccff_tail)
  );


  grid_clb
  grid_clb_7__7_
  (
    .clk_0_N_in(clk_1_wires[151]),
    .prog_clk_0_N_in(prog_clk_1_wires[151]),
    .prog_clk_0_E_out(prog_clk_0_wires[272]),
    .prog_clk_0_S_out(prog_clk_0_wires[271]),
    .config_enable_N_in(config_enableWires[382]),
    .sc_head_S_out(sc_headWires[169]),
    .sc_head_N_in(sc_headWires[168]),
    .reset_E_out(resetWires[168]),
    .reset_W_in(resetWires[167]),
    .Test_en_E_out(Test_enWires[168]),
    .Test_en_W_in(Test_enWires[167]),
    .pReset_N_in(pResetWires[382]),
    .reg_in(reg_out__feedthrough_wires[72]),
    .reg_out(reg_in_feedthrough_wires[71]),
    .cout(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_46_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__65_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_65_ccff_tail)
  );


  grid_clb
  grid_clb_7__8_
  (
    .clk_0_S_in(clk_1_wires[150]),
    .prog_clk_0_S_in(prog_clk_1_wires[150]),
    .prog_clk_0_E_out(prog_clk_0_wires[275]),
    .prog_clk_0_S_out(prog_clk_0_wires[274]),
    .config_enable_N_in(config_enableWires[431]),
    .sc_head_S_out(sc_headWires[167]),
    .sc_head_N_in(sc_headWires[166]),
    .reset_E_out(resetWires[190]),
    .reset_W_in(resetWires[189]),
    .Test_en_E_out(Test_enWires[190]),
    .Test_en_W_in(Test_enWires[189]),
    .pReset_N_in(pResetWires[431]),
    .reg_in(reg_out__feedthrough_wires[73]),
    .reg_out(reg_in_feedthrough_wires[72]),
    .cout(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_47_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__66_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_66_ccff_tail)
  );


  grid_clb
  grid_clb_7__9_
  (
    .clk_0_N_in(clk_1_wires[158]),
    .prog_clk_0_N_in(prog_clk_1_wires[158]),
    .prog_clk_0_E_out(prog_clk_0_wires[278]),
    .prog_clk_0_S_out(prog_clk_0_wires[277]),
    .config_enable_N_in(config_enableWires[480]),
    .sc_head_S_out(sc_headWires[165]),
    .sc_head_N_in(sc_headWires[164]),
    .reset_E_out(resetWires[212]),
    .reset_W_in(resetWires[211]),
    .Test_en_E_out(Test_enWires[212]),
    .Test_en_W_in(Test_enWires[211]),
    .pReset_N_in(pResetWires[480]),
    .reg_in(reg_out__feedthrough_wires[74]),
    .reg_out(reg_in_feedthrough_wires[73]),
    .cout(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_7__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__67_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_67_ccff_tail)
  );


  grid_clb
  grid_clb_7__11_
  (
    .clk_0_N_in(clk_1_wires[165]),
    .prog_clk_0_N_in(prog_clk_1_wires[165]),
    .prog_clk_0_E_out(prog_clk_0_wires[284]),
    .prog_clk_0_S_out(prog_clk_0_wires[283]),
    .config_enable_N_in(config_enableWires[578]),
    .sc_head_S_out(sc_headWires[161]),
    .sc_head_N_in(sc_headWires[160]),
    .reset_E_out(resetWires[256]),
    .reset_W_in(resetWires[255]),
    .Test_en_E_out(Test_enWires[256]),
    .Test_en_W_in(Test_enWires[255]),
    .pReset_N_in(pResetWires[578]),
    .reg_in(reg_out__feedthrough_wires[76]),
    .reg_out(reg_in_feedthrough_wires[75]),
    .cout(grid_clb_7__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_48_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__68_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_68_ccff_tail)
  );


  grid_clb
  grid_clb_7__12_
  (
    .clk_0_S_in(clk_1_wires[164]),
    .prog_clk_0_S_in(prog_clk_1_wires[164]),
    .prog_clk_0_N_out(prog_clk_0_wires[289]),
    .prog_clk_0_E_out(prog_clk_0_wires[287]),
    .prog_clk_0_S_out(prog_clk_0_wires[286]),
    .config_enable_N_in(config_enableWires[621]),
    .sc_head_S_out(sc_headWires[159]),
    .sc_head_N_in(sc_headWires[158]),
    .reset_E_out(resetWires[278]),
    .reset_W_in(resetWires[277]),
    .Test_en_E_out(Test_enWires[278]),
    .Test_en_W_in(Test_enWires[277]),
    .pReset_N_in(pResetWires[621]),
    .reg_out(reg_in_feedthrough_wires[76]),
    .cout(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_7__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__69_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_69_ccff_tail)
  );


  grid_clb
  grid_clb_8__1_
  (
    .clk_0_N_in(clk_1_wires[132]),
    .prog_clk_0_N_in(prog_clk_1_wires[132]),
    .prog_clk_0_E_out(prog_clk_0_wires[292]),
    .prog_clk_0_S_out(prog_clk_0_wires[291]),
    .config_enable_N_in(config_enableWires[92]),
    .sc_head_N_out(sc_headWires[185]),
    .sc_head_S_in(sc_headWires[184]),
    .reset_E_out(resetWires[38]),
    .reset_W_in(resetWires[37]),
    .Test_en_E_out(Test_enWires[38]),
    .Test_en_W_in(Test_enWires[37]),
    .pReset_N_in(pResetWires[92]),
    .reg_in(reg_out__feedthrough_wires[77]),
    .cout(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_49_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__70_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_70_ccff_tail)
  );


  grid_clb
  grid_clb_8__2_
  (
    .clk_0_S_in(clk_1_wires[131]),
    .prog_clk_0_S_in(prog_clk_1_wires[131]),
    .prog_clk_0_E_out(prog_clk_0_wires[295]),
    .prog_clk_0_S_out(prog_clk_0_wires[294]),
    .config_enable_N_in(config_enableWires[141]),
    .sc_head_N_out(sc_headWires[187]),
    .sc_head_S_in(sc_headWires[186]),
    .reset_E_out(resetWires[60]),
    .reset_W_in(resetWires[59]),
    .Test_en_E_out(Test_enWires[60]),
    .Test_en_W_in(Test_enWires[59]),
    .pReset_N_in(pResetWires[141]),
    .reg_in(reg_out__feedthrough_wires[78]),
    .reg_out(reg_in_feedthrough_wires[77]),
    .cout(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__71_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_71_ccff_tail)
  );


  grid_clb
  grid_clb_8__4_
  (
    .clk_0_S_in(clk_1_wires[138]),
    .prog_clk_0_S_in(prog_clk_1_wires[138]),
    .prog_clk_0_E_out(prog_clk_0_wires[301]),
    .prog_clk_0_S_out(prog_clk_0_wires[300]),
    .config_enable_N_in(config_enableWires[239]),
    .sc_head_N_out(sc_headWires[191]),
    .sc_head_S_in(sc_headWires[190]),
    .reset_E_out(resetWires[104]),
    .reset_W_in(resetWires[103]),
    .Test_en_E_out(Test_enWires[104]),
    .Test_en_W_in(Test_enWires[103]),
    .pReset_N_in(pResetWires[239]),
    .reg_in(reg_out__feedthrough_wires[80]),
    .reg_out(reg_in_feedthrough_wires[79]),
    .cout(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_50_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__72_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_72_ccff_tail)
  );


  grid_clb
  grid_clb_8__5_
  (
    .clk_0_N_in(clk_1_wires[146]),
    .prog_clk_0_N_in(prog_clk_1_wires[146]),
    .prog_clk_0_E_out(prog_clk_0_wires[304]),
    .prog_clk_0_S_out(prog_clk_0_wires[303]),
    .config_enable_N_in(config_enableWires[288]),
    .sc_head_N_out(sc_headWires[193]),
    .sc_head_S_in(sc_headWires[192]),
    .reset_E_out(resetWires[126]),
    .reset_W_in(resetWires[125]),
    .Test_en_E_out(Test_enWires[126]),
    .Test_en_W_in(Test_enWires[125]),
    .pReset_N_in(pResetWires[288]),
    .reg_in(reg_out__feedthrough_wires[81]),
    .reg_out(reg_in_feedthrough_wires[80]),
    .cout(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_51_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__73_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_73_ccff_tail)
  );


  grid_clb
  grid_clb_8__6_
  (
    .clk_0_S_in(clk_1_wires[145]),
    .prog_clk_0_S_in(prog_clk_1_wires[145]),
    .prog_clk_0_E_out(prog_clk_0_wires[307]),
    .prog_clk_0_S_out(prog_clk_0_wires[306]),
    .config_enable_N_in(config_enableWires[337]),
    .sc_head_N_out(sc_headWires[195]),
    .sc_head_S_in(sc_headWires[194]),
    .reset_E_out(resetWires[148]),
    .reset_W_in(resetWires[147]),
    .Test_en_E_out(Test_enWires[148]),
    .Test_en_W_in(Test_enWires[147]),
    .pReset_N_in(pResetWires[337]),
    .reg_in(reg_out__feedthrough_wires[82]),
    .reg_out(reg_in_feedthrough_wires[81]),
    .cout(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_52_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__74_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_74_ccff_tail)
  );


  grid_clb
  grid_clb_8__7_
  (
    .clk_0_N_in(clk_1_wires[153]),
    .prog_clk_0_N_in(prog_clk_1_wires[153]),
    .prog_clk_0_E_out(prog_clk_0_wires[310]),
    .prog_clk_0_S_out(prog_clk_0_wires[309]),
    .config_enable_N_in(config_enableWires[386]),
    .sc_head_N_out(sc_headWires[197]),
    .sc_head_S_in(sc_headWires[196]),
    .reset_E_out(resetWires[170]),
    .reset_W_in(resetWires[169]),
    .Test_en_E_out(Test_enWires[170]),
    .Test_en_W_in(Test_enWires[169]),
    .pReset_N_in(pResetWires[386]),
    .reg_in(reg_out__feedthrough_wires[83]),
    .reg_out(reg_in_feedthrough_wires[82]),
    .cout(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_53_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__75_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_75_ccff_tail)
  );


  grid_clb
  grid_clb_8__8_
  (
    .clk_0_S_in(clk_1_wires[152]),
    .prog_clk_0_S_in(prog_clk_1_wires[152]),
    .prog_clk_0_E_out(prog_clk_0_wires[313]),
    .prog_clk_0_S_out(prog_clk_0_wires[312]),
    .config_enable_N_in(config_enableWires[435]),
    .sc_head_N_out(sc_headWires[199]),
    .sc_head_S_in(sc_headWires[198]),
    .reset_E_out(resetWires[192]),
    .reset_W_in(resetWires[191]),
    .Test_en_E_out(Test_enWires[192]),
    .Test_en_W_in(Test_enWires[191]),
    .pReset_N_in(pResetWires[435]),
    .reg_in(reg_out__feedthrough_wires[84]),
    .reg_out(reg_in_feedthrough_wires[83]),
    .cout(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_54_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__76_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_76_ccff_tail)
  );


  grid_clb
  grid_clb_8__9_
  (
    .clk_0_N_in(clk_1_wires[160]),
    .prog_clk_0_N_in(prog_clk_1_wires[160]),
    .prog_clk_0_E_out(prog_clk_0_wires[316]),
    .prog_clk_0_S_out(prog_clk_0_wires[315]),
    .config_enable_N_in(config_enableWires[484]),
    .sc_head_N_out(sc_headWires[201]),
    .sc_head_S_in(sc_headWires[200]),
    .reset_E_out(resetWires[214]),
    .reset_W_in(resetWires[213]),
    .Test_en_E_out(Test_enWires[214]),
    .Test_en_W_in(Test_enWires[213]),
    .pReset_N_in(pResetWires[484]),
    .reg_in(reg_out__feedthrough_wires[85]),
    .reg_out(reg_in_feedthrough_wires[84]),
    .cout(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_8__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__77_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_77_ccff_tail)
  );


  grid_clb
  grid_clb_8__11_
  (
    .clk_0_N_in(clk_1_wires[167]),
    .prog_clk_0_N_in(prog_clk_1_wires[167]),
    .prog_clk_0_E_out(prog_clk_0_wires[322]),
    .prog_clk_0_S_out(prog_clk_0_wires[321]),
    .config_enable_N_in(config_enableWires[582]),
    .sc_head_N_out(sc_headWires[205]),
    .sc_head_S_in(sc_headWires[204]),
    .reset_E_out(resetWires[258]),
    .reset_W_in(resetWires[257]),
    .Test_en_E_out(Test_enWires[258]),
    .Test_en_W_in(Test_enWires[257]),
    .pReset_N_in(pResetWires[582]),
    .reg_in(reg_out__feedthrough_wires[87]),
    .reg_out(reg_in_feedthrough_wires[86]),
    .cout(grid_clb_8__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_55_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__78_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_78_ccff_tail)
  );


  grid_clb
  grid_clb_8__12_
  (
    .clk_0_S_in(clk_1_wires[166]),
    .prog_clk_0_S_in(prog_clk_1_wires[166]),
    .prog_clk_0_N_out(prog_clk_0_wires[327]),
    .prog_clk_0_E_out(prog_clk_0_wires[325]),
    .prog_clk_0_S_out(prog_clk_0_wires[324]),
    .config_enable_N_in(config_enableWires[624]),
    .sc_head_N_out(sc_headWires[207]),
    .sc_head_S_in(sc_headWires[206]),
    .reset_E_out(resetWires[280]),
    .reset_W_in(resetWires[279]),
    .Test_en_E_out(Test_enWires[280]),
    .Test_en_W_in(Test_enWires[279]),
    .pReset_N_in(pResetWires[624]),
    .reg_out(reg_in_feedthrough_wires[87]),
    .cout(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_8__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__79_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_79_ccff_tail)
  );


  grid_clb
  grid_clb_9__1_
  (
    .clk_0_N_in(clk_1_wires[172]),
    .prog_clk_0_N_in(prog_clk_1_wires[172]),
    .prog_clk_0_E_out(prog_clk_0_wires[330]),
    .prog_clk_0_S_out(prog_clk_0_wires[329]),
    .config_enable_N_in(config_enableWires[96]),
    .sc_head_S_out(sc_headWires[233]),
    .sc_head_N_in(sc_headWires[232]),
    .reset_E_out(resetWires[40]),
    .reset_W_in(resetWires[39]),
    .Test_en_E_out(Test_enWires[40]),
    .Test_en_W_in(Test_enWires[39]),
    .pReset_N_in(pResetWires[96]),
    .reg_in(reg_out__feedthrough_wires[88]),
    .cout(grid_clb_9__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_56_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__80_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_80_ccff_tail)
  );


  grid_clb
  grid_clb_9__2_
  (
    .clk_0_S_in(clk_1_wires[171]),
    .prog_clk_0_S_in(prog_clk_1_wires[171]),
    .prog_clk_0_E_out(prog_clk_0_wires[333]),
    .prog_clk_0_S_out(prog_clk_0_wires[332]),
    .config_enable_N_in(config_enableWires[145]),
    .sc_head_S_out(sc_headWires[231]),
    .sc_head_N_in(sc_headWires[230]),
    .reset_E_out(resetWires[62]),
    .reset_W_in(resetWires[61]),
    .Test_en_E_out(Test_enWires[62]),
    .Test_en_W_in(Test_enWires[61]),
    .pReset_N_in(pResetWires[145]),
    .reg_in(reg_out__feedthrough_wires[89]),
    .reg_out(reg_in_feedthrough_wires[88]),
    .cout(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__81_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_81_ccff_tail)
  );


  grid_clb
  grid_clb_9__4_
  (
    .clk_0_S_in(clk_1_wires[178]),
    .prog_clk_0_S_in(prog_clk_1_wires[178]),
    .prog_clk_0_E_out(prog_clk_0_wires[339]),
    .prog_clk_0_S_out(prog_clk_0_wires[338]),
    .config_enable_N_in(config_enableWires[243]),
    .sc_head_S_out(sc_headWires[227]),
    .sc_head_N_in(sc_headWires[226]),
    .reset_E_out(resetWires[106]),
    .reset_W_in(resetWires[105]),
    .Test_en_E_out(Test_enWires[106]),
    .Test_en_W_in(Test_enWires[105]),
    .pReset_N_in(pResetWires[243]),
    .reg_in(reg_out__feedthrough_wires[91]),
    .reg_out(reg_in_feedthrough_wires[90]),
    .cout(grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_57_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__82_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_82_ccff_tail)
  );


  grid_clb
  grid_clb_9__5_
  (
    .clk_0_N_in(clk_1_wires[186]),
    .prog_clk_0_N_in(prog_clk_1_wires[186]),
    .prog_clk_0_E_out(prog_clk_0_wires[342]),
    .prog_clk_0_S_out(prog_clk_0_wires[341]),
    .config_enable_N_in(config_enableWires[292]),
    .sc_head_S_out(sc_headWires[225]),
    .sc_head_N_in(sc_headWires[224]),
    .reset_E_out(resetWires[128]),
    .reset_W_in(resetWires[127]),
    .Test_en_E_out(Test_enWires[128]),
    .Test_en_W_in(Test_enWires[127]),
    .pReset_N_in(pResetWires[292]),
    .reg_in(reg_out__feedthrough_wires[92]),
    .reg_out(reg_in_feedthrough_wires[91]),
    .cout(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_58_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__83_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_83_ccff_tail)
  );


  grid_clb
  grid_clb_9__6_
  (
    .clk_0_S_in(clk_1_wires[185]),
    .prog_clk_0_S_in(prog_clk_1_wires[185]),
    .prog_clk_0_E_out(prog_clk_0_wires[345]),
    .prog_clk_0_S_out(prog_clk_0_wires[344]),
    .config_enable_N_in(config_enableWires[341]),
    .sc_head_S_out(sc_headWires[223]),
    .sc_head_N_in(sc_headWires[222]),
    .reset_E_out(resetWires[150]),
    .reset_W_in(resetWires[149]),
    .Test_en_E_out(Test_enWires[150]),
    .Test_en_W_in(Test_enWires[149]),
    .pReset_N_in(pResetWires[341]),
    .reg_in(reg_out__feedthrough_wires[93]),
    .reg_out(reg_in_feedthrough_wires[92]),
    .cout(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_59_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__84_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_84_ccff_tail)
  );


  grid_clb
  grid_clb_9__7_
  (
    .clk_0_N_in(clk_1_wires[193]),
    .prog_clk_0_N_in(prog_clk_1_wires[193]),
    .prog_clk_0_E_out(prog_clk_0_wires[348]),
    .prog_clk_0_S_out(prog_clk_0_wires[347]),
    .config_enable_N_in(config_enableWires[390]),
    .sc_head_S_out(sc_headWires[221]),
    .sc_head_N_in(sc_headWires[220]),
    .reset_E_out(resetWires[172]),
    .reset_W_in(resetWires[171]),
    .Test_en_E_out(Test_enWires[172]),
    .Test_en_W_in(Test_enWires[171]),
    .pReset_N_in(pResetWires[390]),
    .reg_in(reg_out__feedthrough_wires[94]),
    .reg_out(reg_in_feedthrough_wires[93]),
    .cout(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_60_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__85_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_85_ccff_tail)
  );


  grid_clb
  grid_clb_9__8_
  (
    .clk_0_S_in(clk_1_wires[192]),
    .prog_clk_0_S_in(prog_clk_1_wires[192]),
    .prog_clk_0_E_out(prog_clk_0_wires[351]),
    .prog_clk_0_S_out(prog_clk_0_wires[350]),
    .config_enable_N_in(config_enableWires[439]),
    .sc_head_S_out(sc_headWires[219]),
    .sc_head_N_in(sc_headWires[218]),
    .reset_E_out(resetWires[194]),
    .reset_W_in(resetWires[193]),
    .Test_en_E_out(Test_enWires[194]),
    .Test_en_W_in(Test_enWires[193]),
    .pReset_N_in(pResetWires[439]),
    .reg_in(reg_out__feedthrough_wires[95]),
    .reg_out(reg_in_feedthrough_wires[94]),
    .cout(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_61_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__86_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_86_ccff_tail)
  );


  grid_clb
  grid_clb_9__9_
  (
    .clk_0_N_in(clk_1_wires[200]),
    .prog_clk_0_N_in(prog_clk_1_wires[200]),
    .prog_clk_0_E_out(prog_clk_0_wires[354]),
    .prog_clk_0_S_out(prog_clk_0_wires[353]),
    .config_enable_N_in(config_enableWires[488]),
    .sc_head_S_out(sc_headWires[217]),
    .sc_head_N_in(sc_headWires[216]),
    .reset_E_out(resetWires[216]),
    .reset_W_in(resetWires[215]),
    .Test_en_E_out(Test_enWires[216]),
    .Test_en_W_in(Test_enWires[215]),
    .pReset_N_in(pResetWires[488]),
    .reg_in(reg_out__feedthrough_wires[96]),
    .reg_out(reg_in_feedthrough_wires[95]),
    .cout(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_9__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__87_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_87_ccff_tail)
  );


  grid_clb
  grid_clb_9__11_
  (
    .clk_0_N_in(clk_1_wires[207]),
    .prog_clk_0_N_in(prog_clk_1_wires[207]),
    .prog_clk_0_E_out(prog_clk_0_wires[360]),
    .prog_clk_0_S_out(prog_clk_0_wires[359]),
    .config_enable_N_in(config_enableWires[586]),
    .sc_head_S_out(sc_headWires[213]),
    .sc_head_N_in(sc_headWires[212]),
    .reset_E_out(resetWires[260]),
    .reset_W_in(resetWires[259]),
    .Test_en_E_out(Test_enWires[260]),
    .Test_en_W_in(Test_enWires[259]),
    .pReset_N_in(pResetWires[586]),
    .reg_in(reg_out__feedthrough_wires[98]),
    .reg_out(reg_in_feedthrough_wires[97]),
    .cout(grid_clb_9__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_62_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__88_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_88_ccff_tail)
  );


  grid_clb
  grid_clb_9__12_
  (
    .clk_0_S_in(clk_1_wires[206]),
    .prog_clk_0_S_in(prog_clk_1_wires[206]),
    .prog_clk_0_N_out(prog_clk_0_wires[365]),
    .prog_clk_0_E_out(prog_clk_0_wires[363]),
    .prog_clk_0_S_out(prog_clk_0_wires[362]),
    .config_enable_N_in(config_enableWires[627]),
    .sc_head_S_out(sc_headWires[211]),
    .sc_head_N_in(sc_headWires[210]),
    .reset_E_out(resetWires[282]),
    .reset_W_in(resetWires[281]),
    .Test_en_E_out(Test_enWires[282]),
    .Test_en_W_in(Test_enWires[281]),
    .pReset_N_in(pResetWires[627]),
    .reg_out(reg_in_feedthrough_wires[98]),
    .cout(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_9__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__89_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_89_ccff_tail)
  );


  grid_clb
  grid_clb_10__1_
  (
    .clk_0_N_in(clk_1_wires[174]),
    .prog_clk_0_N_in(prog_clk_1_wires[174]),
    .prog_clk_0_E_out(prog_clk_0_wires[368]),
    .prog_clk_0_S_out(prog_clk_0_wires[367]),
    .config_enable_N_in(config_enableWires[100]),
    .sc_head_N_out(sc_headWires[237]),
    .sc_head_S_in(sc_headWires[236]),
    .reset_E_out(resetWires[42]),
    .reset_W_in(resetWires[41]),
    .Test_en_E_out(Test_enWires[42]),
    .Test_en_W_in(Test_enWires[41]),
    .pReset_N_in(pResetWires[100]),
    .reg_in(reg_out__feedthrough_wires[99]),
    .cout(grid_clb_10__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_63_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__90_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_90_ccff_tail)
  );


  grid_clb
  grid_clb_10__2_
  (
    .clk_0_S_in(clk_1_wires[173]),
    .prog_clk_0_S_in(prog_clk_1_wires[173]),
    .prog_clk_0_E_out(prog_clk_0_wires[371]),
    .prog_clk_0_S_out(prog_clk_0_wires[370]),
    .config_enable_N_in(config_enableWires[149]),
    .sc_head_N_out(sc_headWires[239]),
    .sc_head_S_in(sc_headWires[238]),
    .reset_E_out(resetWires[64]),
    .reset_W_in(resetWires[63]),
    .Test_en_E_out(Test_enWires[64]),
    .Test_en_W_in(Test_enWires[63]),
    .pReset_N_in(pResetWires[149]),
    .reg_in(reg_out__feedthrough_wires[100]),
    .reg_out(reg_in_feedthrough_wires[99]),
    .cout(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_10__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__91_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_91_ccff_tail)
  );


  grid_clb
  grid_clb_10__4_
  (
    .clk_0_S_in(clk_1_wires[180]),
    .prog_clk_0_S_in(prog_clk_1_wires[180]),
    .prog_clk_0_E_out(prog_clk_0_wires[377]),
    .prog_clk_0_S_out(prog_clk_0_wires[376]),
    .config_enable_N_in(config_enableWires[247]),
    .sc_head_N_out(sc_headWires[243]),
    .sc_head_S_in(sc_headWires[242]),
    .reset_E_out(resetWires[108]),
    .reset_W_in(resetWires[107]),
    .Test_en_E_out(Test_enWires[108]),
    .Test_en_W_in(Test_enWires[107]),
    .pReset_N_in(pResetWires[247]),
    .reg_in(reg_out__feedthrough_wires[102]),
    .reg_out(reg_in_feedthrough_wires[101]),
    .cout(grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_64_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__92_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_92_ccff_tail)
  );


  grid_clb
  grid_clb_10__5_
  (
    .clk_0_N_in(clk_1_wires[188]),
    .prog_clk_0_N_in(prog_clk_1_wires[188]),
    .prog_clk_0_E_out(prog_clk_0_wires[380]),
    .prog_clk_0_S_out(prog_clk_0_wires[379]),
    .config_enable_N_in(config_enableWires[296]),
    .sc_head_N_out(sc_headWires[245]),
    .sc_head_S_in(sc_headWires[244]),
    .reset_E_out(resetWires[130]),
    .reset_W_in(resetWires[129]),
    .Test_en_E_out(Test_enWires[130]),
    .Test_en_W_in(Test_enWires[129]),
    .pReset_N_in(pResetWires[296]),
    .reg_in(reg_out__feedthrough_wires[103]),
    .reg_out(reg_in_feedthrough_wires[102]),
    .cout(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_65_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__93_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_93_ccff_tail)
  );


  grid_clb
  grid_clb_10__6_
  (
    .clk_0_S_in(clk_1_wires[187]),
    .prog_clk_0_S_in(prog_clk_1_wires[187]),
    .prog_clk_0_E_out(prog_clk_0_wires[383]),
    .prog_clk_0_S_out(prog_clk_0_wires[382]),
    .config_enable_N_in(config_enableWires[345]),
    .sc_head_N_out(sc_headWires[247]),
    .sc_head_S_in(sc_headWires[246]),
    .reset_E_out(resetWires[152]),
    .reset_W_in(resetWires[151]),
    .Test_en_E_out(Test_enWires[152]),
    .Test_en_W_in(Test_enWires[151]),
    .pReset_N_in(pResetWires[345]),
    .reg_in(reg_out__feedthrough_wires[104]),
    .reg_out(reg_in_feedthrough_wires[103]),
    .cout(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_66_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__94_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_94_ccff_tail)
  );


  grid_clb
  grid_clb_10__7_
  (
    .clk_0_N_in(clk_1_wires[195]),
    .prog_clk_0_N_in(prog_clk_1_wires[195]),
    .prog_clk_0_E_out(prog_clk_0_wires[386]),
    .prog_clk_0_S_out(prog_clk_0_wires[385]),
    .config_enable_N_in(config_enableWires[394]),
    .sc_head_N_out(sc_headWires[249]),
    .sc_head_S_in(sc_headWires[248]),
    .reset_E_out(resetWires[174]),
    .reset_W_in(resetWires[173]),
    .Test_en_E_out(Test_enWires[174]),
    .Test_en_W_in(Test_enWires[173]),
    .pReset_N_in(pResetWires[394]),
    .reg_in(reg_out__feedthrough_wires[105]),
    .reg_out(reg_in_feedthrough_wires[104]),
    .cout(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_67_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__95_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_95_ccff_tail)
  );


  grid_clb
  grid_clb_10__8_
  (
    .clk_0_S_in(clk_1_wires[194]),
    .prog_clk_0_S_in(prog_clk_1_wires[194]),
    .prog_clk_0_E_out(prog_clk_0_wires[389]),
    .prog_clk_0_S_out(prog_clk_0_wires[388]),
    .config_enable_N_in(config_enableWires[443]),
    .sc_head_N_out(sc_headWires[251]),
    .sc_head_S_in(sc_headWires[250]),
    .reset_E_out(resetWires[196]),
    .reset_W_in(resetWires[195]),
    .Test_en_E_out(Test_enWires[196]),
    .Test_en_W_in(Test_enWires[195]),
    .pReset_N_in(pResetWires[443]),
    .reg_in(reg_out__feedthrough_wires[106]),
    .reg_out(reg_in_feedthrough_wires[105]),
    .cout(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_68_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__96_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_96_ccff_tail)
  );


  grid_clb
  grid_clb_10__9_
  (
    .clk_0_N_in(clk_1_wires[202]),
    .prog_clk_0_N_in(prog_clk_1_wires[202]),
    .prog_clk_0_E_out(prog_clk_0_wires[392]),
    .prog_clk_0_S_out(prog_clk_0_wires[391]),
    .config_enable_N_in(config_enableWires[492]),
    .sc_head_N_out(sc_headWires[253]),
    .sc_head_S_in(sc_headWires[252]),
    .reset_E_out(resetWires[218]),
    .reset_W_in(resetWires[217]),
    .Test_en_E_out(Test_enWires[218]),
    .Test_en_W_in(Test_enWires[217]),
    .pReset_N_in(pResetWires[492]),
    .reg_in(reg_out__feedthrough_wires[107]),
    .reg_out(reg_in_feedthrough_wires[106]),
    .cout(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_10__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__97_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_97_ccff_tail)
  );


  grid_clb
  grid_clb_10__11_
  (
    .clk_0_N_in(clk_1_wires[209]),
    .prog_clk_0_N_in(prog_clk_1_wires[209]),
    .prog_clk_0_E_out(prog_clk_0_wires[398]),
    .prog_clk_0_S_out(prog_clk_0_wires[397]),
    .config_enable_N_in(config_enableWires[590]),
    .sc_head_N_out(sc_headWires[257]),
    .sc_head_S_in(sc_headWires[256]),
    .reset_E_out(resetWires[262]),
    .reset_W_in(resetWires[261]),
    .Test_en_E_out(Test_enWires[262]),
    .Test_en_W_in(Test_enWires[261]),
    .pReset_N_in(pResetWires[590]),
    .reg_in(reg_out__feedthrough_wires[109]),
    .reg_out(reg_in_feedthrough_wires[108]),
    .cout(grid_clb_10__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_69_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__98_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_98_ccff_tail)
  );


  grid_clb
  grid_clb_10__12_
  (
    .clk_0_S_in(clk_1_wires[208]),
    .prog_clk_0_S_in(prog_clk_1_wires[208]),
    .prog_clk_0_N_out(prog_clk_0_wires[403]),
    .prog_clk_0_E_out(prog_clk_0_wires[401]),
    .prog_clk_0_S_out(prog_clk_0_wires[400]),
    .config_enable_N_in(config_enableWires[630]),
    .sc_head_N_out(sc_headWires[259]),
    .sc_head_S_in(sc_headWires[258]),
    .reset_E_out(resetWires[284]),
    .reset_W_in(resetWires[283]),
    .Test_en_E_out(Test_enWires[284]),
    .Test_en_W_in(Test_enWires[283]),
    .pReset_N_in(pResetWires[630]),
    .reg_out(reg_in_feedthrough_wires[109]),
    .cout(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_10__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__99_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_99_ccff_tail)
  );


  grid_clb
  grid_clb_11__1_
  (
    .clk_0_N_in(clk_1_wires[214]),
    .prog_clk_0_N_in(prog_clk_1_wires[214]),
    .prog_clk_0_E_out(prog_clk_0_wires[406]),
    .prog_clk_0_S_out(prog_clk_0_wires[405]),
    .config_enable_N_in(config_enableWires[104]),
    .sc_head_S_out(sc_headWires[285]),
    .sc_head_N_in(sc_headWires[284]),
    .reset_E_out(resetWires[44]),
    .reset_W_in(resetWires[43]),
    .Test_en_E_out(Test_enWires[44]),
    .Test_en_W_in(Test_enWires[43]),
    .pReset_N_in(pResetWires[104]),
    .reg_in(reg_out__feedthrough_wires[110]),
    .cout(grid_clb_11__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_70_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__100_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_100_ccff_tail)
  );


  grid_clb
  grid_clb_11__2_
  (
    .clk_0_S_in(clk_1_wires[213]),
    .prog_clk_0_S_in(prog_clk_1_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[409]),
    .prog_clk_0_S_out(prog_clk_0_wires[408]),
    .config_enable_N_in(config_enableWires[153]),
    .sc_head_S_out(sc_headWires[283]),
    .sc_head_N_in(sc_headWires[282]),
    .reset_E_out(resetWires[66]),
    .reset_W_in(resetWires[65]),
    .Test_en_E_out(Test_enWires[66]),
    .Test_en_W_in(Test_enWires[65]),
    .pReset_N_in(pResetWires[153]),
    .reg_in(reg_out__feedthrough_wires[111]),
    .reg_out(reg_in_feedthrough_wires[110]),
    .cout(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_11__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__101_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_101_ccff_tail)
  );


  grid_clb
  grid_clb_11__4_
  (
    .clk_0_S_in(clk_1_wires[220]),
    .prog_clk_0_S_in(prog_clk_1_wires[220]),
    .prog_clk_0_E_out(prog_clk_0_wires[415]),
    .prog_clk_0_S_out(prog_clk_0_wires[414]),
    .config_enable_N_in(config_enableWires[251]),
    .sc_head_S_out(sc_headWires[279]),
    .sc_head_N_in(sc_headWires[278]),
    .reset_E_out(resetWires[110]),
    .reset_W_in(resetWires[109]),
    .Test_en_E_out(Test_enWires[110]),
    .Test_en_W_in(Test_enWires[109]),
    .pReset_N_in(pResetWires[251]),
    .reg_in(reg_out__feedthrough_wires[113]),
    .reg_out(reg_in_feedthrough_wires[112]),
    .cout(grid_clb_11__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_71_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__102_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_102_ccff_tail)
  );


  grid_clb
  grid_clb_11__5_
  (
    .clk_0_N_in(clk_1_wires[228]),
    .prog_clk_0_N_in(prog_clk_1_wires[228]),
    .prog_clk_0_E_out(prog_clk_0_wires[418]),
    .prog_clk_0_S_out(prog_clk_0_wires[417]),
    .config_enable_N_in(config_enableWires[300]),
    .sc_head_S_out(sc_headWires[277]),
    .sc_head_N_in(sc_headWires[276]),
    .reset_E_out(resetWires[132]),
    .reset_W_in(resetWires[131]),
    .Test_en_E_out(Test_enWires[132]),
    .Test_en_W_in(Test_enWires[131]),
    .pReset_N_in(pResetWires[300]),
    .reg_in(reg_out__feedthrough_wires[114]),
    .reg_out(reg_in_feedthrough_wires[113]),
    .cout(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_72_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__103_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_103_ccff_tail)
  );


  grid_clb
  grid_clb_11__6_
  (
    .clk_0_S_in(clk_1_wires[227]),
    .prog_clk_0_S_in(prog_clk_1_wires[227]),
    .prog_clk_0_E_out(prog_clk_0_wires[421]),
    .prog_clk_0_S_out(prog_clk_0_wires[420]),
    .config_enable_N_in(config_enableWires[349]),
    .sc_head_S_out(sc_headWires[275]),
    .sc_head_N_in(sc_headWires[274]),
    .reset_E_out(resetWires[154]),
    .reset_W_in(resetWires[153]),
    .Test_en_E_out(Test_enWires[154]),
    .Test_en_W_in(Test_enWires[153]),
    .pReset_N_in(pResetWires[349]),
    .reg_in(reg_out__feedthrough_wires[115]),
    .reg_out(reg_in_feedthrough_wires[114]),
    .cout(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_73_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__104_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_104_ccff_tail)
  );


  grid_clb
  grid_clb_11__7_
  (
    .clk_0_N_in(clk_1_wires[235]),
    .prog_clk_0_N_in(prog_clk_1_wires[235]),
    .prog_clk_0_E_out(prog_clk_0_wires[424]),
    .prog_clk_0_S_out(prog_clk_0_wires[423]),
    .config_enable_N_in(config_enableWires[398]),
    .sc_head_S_out(sc_headWires[273]),
    .sc_head_N_in(sc_headWires[272]),
    .reset_E_out(resetWires[176]),
    .reset_W_in(resetWires[175]),
    .Test_en_E_out(Test_enWires[176]),
    .Test_en_W_in(Test_enWires[175]),
    .pReset_N_in(pResetWires[398]),
    .reg_in(reg_out__feedthrough_wires[116]),
    .reg_out(reg_in_feedthrough_wires[115]),
    .cout(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_74_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__105_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_105_ccff_tail)
  );


  grid_clb
  grid_clb_11__8_
  (
    .clk_0_S_in(clk_1_wires[234]),
    .prog_clk_0_S_in(prog_clk_1_wires[234]),
    .prog_clk_0_E_out(prog_clk_0_wires[427]),
    .prog_clk_0_S_out(prog_clk_0_wires[426]),
    .config_enable_N_in(config_enableWires[447]),
    .sc_head_S_out(sc_headWires[271]),
    .sc_head_N_in(sc_headWires[270]),
    .reset_E_out(resetWires[198]),
    .reset_W_in(resetWires[197]),
    .Test_en_E_out(Test_enWires[198]),
    .Test_en_W_in(Test_enWires[197]),
    .pReset_N_in(pResetWires[447]),
    .reg_in(reg_out__feedthrough_wires[117]),
    .reg_out(reg_in_feedthrough_wires[116]),
    .cout(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_75_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__106_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_106_ccff_tail)
  );


  grid_clb
  grid_clb_11__9_
  (
    .clk_0_N_in(clk_1_wires[242]),
    .prog_clk_0_N_in(prog_clk_1_wires[242]),
    .prog_clk_0_E_out(prog_clk_0_wires[430]),
    .prog_clk_0_S_out(prog_clk_0_wires[429]),
    .config_enable_N_in(config_enableWires[496]),
    .sc_head_S_out(sc_headWires[269]),
    .sc_head_N_in(sc_headWires[268]),
    .reset_E_out(resetWires[220]),
    .reset_W_in(resetWires[219]),
    .Test_en_E_out(Test_enWires[220]),
    .Test_en_W_in(Test_enWires[219]),
    .pReset_N_in(pResetWires[496]),
    .reg_in(reg_out__feedthrough_wires[118]),
    .reg_out(reg_in_feedthrough_wires[117]),
    .cout(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_11__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__107_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_107_ccff_tail)
  );


  grid_clb
  grid_clb_11__11_
  (
    .clk_0_N_in(clk_1_wires[249]),
    .prog_clk_0_N_in(prog_clk_1_wires[249]),
    .prog_clk_0_E_out(prog_clk_0_wires[436]),
    .prog_clk_0_S_out(prog_clk_0_wires[435]),
    .config_enable_N_in(config_enableWires[594]),
    .sc_head_S_out(sc_headWires[265]),
    .sc_head_N_in(sc_headWires[264]),
    .reset_E_out(resetWires[264]),
    .reset_W_in(resetWires[263]),
    .Test_en_E_out(Test_enWires[264]),
    .Test_en_W_in(Test_enWires[263]),
    .pReset_N_in(pResetWires[594]),
    .reg_in(reg_out__feedthrough_wires[120]),
    .reg_out(reg_in_feedthrough_wires[119]),
    .cout(grid_clb_11__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_76_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__108_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_108_ccff_tail)
  );


  grid_clb
  grid_clb_11__12_
  (
    .clk_0_S_in(clk_1_wires[248]),
    .prog_clk_0_S_in(prog_clk_1_wires[248]),
    .prog_clk_0_N_out(prog_clk_0_wires[441]),
    .prog_clk_0_E_out(prog_clk_0_wires[439]),
    .prog_clk_0_S_out(prog_clk_0_wires[438]),
    .config_enable_N_in(config_enableWires[633]),
    .sc_head_S_out(sc_headWires[263]),
    .sc_head_N_in(sc_headWires[262]),
    .reset_E_out(resetWires[286]),
    .reset_W_in(resetWires[285]),
    .Test_en_E_out(Test_enWires[286]),
    .Test_en_W_in(Test_enWires[285]),
    .pReset_N_in(pResetWires[633]),
    .reg_out(reg_in_feedthrough_wires[120]),
    .cout(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_11__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(cby_1__1__109_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_109_ccff_tail)
  );


  grid_clb
  grid_clb_12__1_
  (
    .clk_0_N_in(clk_1_wires[216]),
    .prog_clk_0_N_in(prog_clk_1_wires[216]),
    .prog_clk_0_E_out(prog_clk_0_wires[444]),
    .prog_clk_0_S_out(prog_clk_0_wires[443]),
    .config_enable_N_in(config_enableWires[108]),
    .sc_head_N_out(sc_headWires[289]),
    .sc_head_S_in(sc_headWires[288]),
    .reset_W_in(resetWires[45]),
    .Test_en_W_in(Test_enWires[45]),
    .pReset_N_in(pResetWires[108]),
    .reg_in(reg_out__feedthrough_wires[121]),
    .cout(grid_clb_12__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_77_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_11_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_110_ccff_tail)
  );


  grid_clb
  grid_clb_12__2_
  (
    .clk_0_S_in(clk_1_wires[215]),
    .prog_clk_0_S_in(prog_clk_1_wires[215]),
    .prog_clk_0_E_out(prog_clk_0_wires[447]),
    .prog_clk_0_S_out(prog_clk_0_wires[446]),
    .config_enable_N_in(config_enableWires[157]),
    .sc_head_N_out(sc_headWires[291]),
    .sc_head_S_in(sc_headWires[290]),
    .reset_W_in(resetWires[67]),
    .Test_en_W_in(Test_enWires[67]),
    .pReset_N_in(pResetWires[157]),
    .reg_in(reg_out__feedthrough_wires[122]),
    .reg_out(reg_in_feedthrough_wires[121]),
    .cout(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_12__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_10_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_111_ccff_tail)
  );


  grid_clb
  grid_clb_12__4_
  (
    .clk_0_S_in(clk_1_wires[222]),
    .prog_clk_0_S_in(prog_clk_1_wires[222]),
    .prog_clk_0_E_out(prog_clk_0_wires[453]),
    .prog_clk_0_S_out(prog_clk_0_wires[452]),
    .config_enable_N_in(config_enableWires[255]),
    .sc_head_N_out(sc_headWires[295]),
    .sc_head_S_in(sc_headWires[294]),
    .reset_W_in(resetWires[111]),
    .Test_en_W_in(Test_enWires[111]),
    .pReset_N_in(pResetWires[255]),
    .reg_in(reg_out__feedthrough_wires[124]),
    .reg_out(reg_in_feedthrough_wires[123]),
    .cout(grid_clb_12__4__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_78_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_112_ccff_tail)
  );


  grid_clb
  grid_clb_12__5_
  (
    .clk_0_N_in(clk_1_wires[230]),
    .prog_clk_0_N_in(prog_clk_1_wires[230]),
    .prog_clk_0_E_out(prog_clk_0_wires[456]),
    .prog_clk_0_S_out(prog_clk_0_wires[455]),
    .config_enable_N_in(config_enableWires[304]),
    .sc_head_N_out(sc_headWires[297]),
    .sc_head_S_in(sc_headWires[296]),
    .reset_W_in(resetWires[133]),
    .Test_en_W_in(Test_enWires[133]),
    .pReset_N_in(pResetWires[304]),
    .reg_in(reg_out__feedthrough_wires[125]),
    .reg_out(reg_in_feedthrough_wires[124]),
    .cout(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_79_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_113_ccff_tail)
  );


  grid_clb
  grid_clb_12__6_
  (
    .clk_0_S_in(clk_1_wires[229]),
    .prog_clk_0_S_in(prog_clk_1_wires[229]),
    .prog_clk_0_E_out(prog_clk_0_wires[459]),
    .prog_clk_0_S_out(prog_clk_0_wires[458]),
    .config_enable_N_in(config_enableWires[353]),
    .sc_head_N_out(sc_headWires[299]),
    .sc_head_S_in(sc_headWires[298]),
    .reset_W_in(resetWires[155]),
    .Test_en_W_in(Test_enWires[155]),
    .pReset_N_in(pResetWires[353]),
    .reg_in(reg_out__feedthrough_wires[126]),
    .reg_out(reg_in_feedthrough_wires[125]),
    .cout(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_80_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_114_ccff_tail)
  );


  grid_clb
  grid_clb_12__7_
  (
    .clk_0_N_in(clk_1_wires[237]),
    .prog_clk_0_N_in(prog_clk_1_wires[237]),
    .prog_clk_0_E_out(prog_clk_0_wires[462]),
    .prog_clk_0_S_out(prog_clk_0_wires[461]),
    .config_enable_N_in(config_enableWires[402]),
    .sc_head_N_out(sc_headWires[301]),
    .sc_head_S_in(sc_headWires[300]),
    .reset_W_in(resetWires[177]),
    .Test_en_W_in(Test_enWires[177]),
    .pReset_N_in(pResetWires[402]),
    .reg_in(reg_out__feedthrough_wires[127]),
    .reg_out(reg_in_feedthrough_wires[126]),
    .cout(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_81_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_115_ccff_tail)
  );


  grid_clb
  grid_clb_12__8_
  (
    .clk_0_S_in(clk_1_wires[236]),
    .prog_clk_0_S_in(prog_clk_1_wires[236]),
    .prog_clk_0_E_out(prog_clk_0_wires[465]),
    .prog_clk_0_S_out(prog_clk_0_wires[464]),
    .config_enable_N_in(config_enableWires[451]),
    .sc_head_N_out(sc_headWires[303]),
    .sc_head_S_in(sc_headWires[302]),
    .reset_W_in(resetWires[199]),
    .Test_en_W_in(Test_enWires[199]),
    .pReset_N_in(pResetWires[451]),
    .reg_in(reg_out__feedthrough_wires[128]),
    .reg_out(reg_in_feedthrough_wires[127]),
    .cout(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_82_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_116_ccff_tail)
  );


  grid_clb
  grid_clb_12__9_
  (
    .clk_0_N_in(clk_1_wires[244]),
    .prog_clk_0_N_in(prog_clk_1_wires[244]),
    .prog_clk_0_E_out(prog_clk_0_wires[468]),
    .prog_clk_0_S_out(prog_clk_0_wires[467]),
    .config_enable_N_in(config_enableWires[500]),
    .sc_head_N_out(sc_headWires[305]),
    .sc_head_S_in(sc_headWires[304]),
    .reset_W_in(resetWires[221]),
    .Test_en_W_in(Test_enWires[221]),
    .pReset_N_in(pResetWires[500]),
    .reg_in(reg_out__feedthrough_wires[129]),
    .reg_out(reg_in_feedthrough_wires[128]),
    .cout(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_12__9__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_117_ccff_tail)
  );


  grid_clb
  grid_clb_12__11_
  (
    .clk_0_N_in(clk_1_wires[251]),
    .prog_clk_0_N_in(prog_clk_1_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[474]),
    .prog_clk_0_S_out(prog_clk_0_wires[473]),
    .config_enable_N_in(config_enableWires[598]),
    .sc_head_N_out(sc_headWires[309]),
    .sc_head_S_in(sc_headWires[308]),
    .reset_W_in(resetWires[265]),
    .Test_en_W_in(Test_enWires[265]),
    .pReset_N_in(pResetWires[598]),
    .reg_in(reg_out__feedthrough_wires[131]),
    .reg_out(reg_in_feedthrough_wires[130]),
    .cout(grid_clb_12__11__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(direct_interc_83_out),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_118_ccff_tail)
  );


  grid_clb
  grid_clb_12__12_
  (
    .clk_0_S_in(clk_1_wires[250]),
    .prog_clk_0_S_in(prog_clk_1_wires[250]),
    .prog_clk_0_N_out(prog_clk_0_wires[479]),
    .prog_clk_0_E_out(prog_clk_0_wires[477]),
    .prog_clk_0_S_out(prog_clk_0_wires[476]),
    .config_enable_N_in(config_enableWires[636]),
    .sc_head_N_out(sc_headWires[311]),
    .sc_head_S_in(sc_headWires[310]),
    .reset_W_in(resetWires[287]),
    .Test_en_W_in(Test_enWires[287]),
    .pReset_N_in(pResetWires[636]),
    .reg_out(reg_in_feedthrough_wires[131]),
    .cout(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .cin(grid_clb_12__12__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
    .top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__12__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .right_width_0_height_0_subtile_0__pin_I_9_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .right_width_0_height_0_subtile_0__pin_I_10_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .right_width_0_height_0_subtile_0__pin_I_11_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .right_width_0_height_0_subtile_0__pin_I_12_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .right_width_0_height_0_subtile_0__pin_I_13_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .right_width_0_height_0_subtile_0__pin_I_14_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .right_width_0_height_0_subtile_0__pin_I_15_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .right_width_0_height_0_subtile_0__pin_I_16_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .right_width_0_height_0_subtile_0__pin_I_17_(cby_12__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_head(grid_io_right_right_0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .right_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .right_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .right_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .right_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .ccff_tail(grid_clb_119_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_1__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__0_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__0_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__0_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__0_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[114]),
    .cby_config_enable_S_in_in_1(config_enableWires[114]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[13]),
    .grid_clb_pReset_N_in_in_2(pResetWires[166]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[69]),
    .grid_clb_reset_E_in_in_2(resetWires[69]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[32]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[33]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[166]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[69]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[70]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[13]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[13]),
    .grid_clb_pReset_N_in_in_1(pResetWires[161]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[20]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[21]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[161]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[11]),
    .grid_clb_prog_clk_0_W_out_out_1(prog_clk_0_wires[14]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[11]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[11]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__0_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_0_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_1__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__1_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__1_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__1_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__1_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[457]),
    .cby_config_enable_S_in_in_1(config_enableWires[457]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[48]),
    .grid_clb_pReset_N_in_in_2(pResetWires[509]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[223]),
    .grid_clb_reset_E_in_in_2(resetWires[223]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[46]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[47]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[509]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[90]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[91]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[33]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[33]),
    .grid_clb_pReset_N_in_in_1(pResetWires[504]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[6]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[7]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[504]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[46]),
    .grid_clb_prog_clk_0_W_out_out_1(prog_clk_0_wires[49]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[31]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[31]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__1_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_1_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_3__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__2_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__2_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__2_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__2_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[122]),
    .cby_config_enable_S_in_in_1(config_enableWires[122]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[109]),
    .grid_clb_pReset_N_in_in_2(pResetWires[174]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[73]),
    .grid_clb_reset_E_in_in_2(resetWires[73]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[84]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[85]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[174]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[145]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[146]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[55]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[55]),
    .grid_clb_pReset_N_in_in_1(pResetWires[170]),
    .grid_clb_Test_en_W_out_out_1(Test_enWires[72]),
    .grid_clb_reset_W_out_out_1(resetWires[72]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[72]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[73]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[170]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[107]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[53]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[53]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_2_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_3__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__3_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__3_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__3_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__3_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[465]),
    .cby_config_enable_S_in_in_1(config_enableWires[465]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[130]),
    .grid_clb_pReset_N_in_in_2(pResetWires[517]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[227]),
    .grid_clb_reset_E_in_in_2(resetWires[227]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[98]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[99]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[517]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[166]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[167]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[75]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[75]),
    .grid_clb_pReset_N_in_in_1(pResetWires[513]),
    .grid_clb_Test_en_W_out_out_1(Test_enWires[226]),
    .grid_clb_reset_W_out_out_1(resetWires[226]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[58]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[59]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[513]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[128]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[73]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[73]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__3_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_3_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_5__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__4_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__4_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__4_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__4_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[130]),
    .cby_config_enable_S_in_in_1(config_enableWires[130]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[185]),
    .grid_clb_pReset_N_in_in_2(pResetWires[182]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[77]),
    .grid_clb_reset_E_in_in_2(resetWires[77]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[136]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[137]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[182]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[221]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[222]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[97]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[97]),
    .grid_clb_pReset_N_in_in_1(pResetWires[178]),
    .grid_clb_Test_en_W_out_out_1(Test_enWires[76]),
    .grid_clb_reset_W_out_out_1(resetWires[76]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[124]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[125]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[178]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[183]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[95]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[95]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__4_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_4_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_5__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__5_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__5_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__5_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__5_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[473]),
    .cby_config_enable_S_in_in_1(config_enableWires[473]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[206]),
    .grid_clb_pReset_N_in_in_2(pResetWires[525]),
    .grid_clb_Test_en_E_in_in_2(Test_enWires[231]),
    .grid_clb_reset_E_in_in_2(resetWires[231]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[150]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[151]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[525]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[242]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[243]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[117]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[117]),
    .grid_clb_pReset_N_in_in_1(pResetWires[521]),
    .grid_clb_Test_en_W_out_out_1(Test_enWires[230]),
    .grid_clb_reset_W_out_out_1(resetWires[230]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[110]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[111]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[521]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[204]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[115]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[115]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__5_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_5_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_7__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__6_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__6_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__6_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__6_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[138]),
    .cby_config_enable_S_in_in_1(config_enableWires[138]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[261]),
    .grid_clb_pReset_N_in_in_2(pResetWires[190]),
    .grid_clb_Test_en_E_out_out_2(Test_enWires[82]),
    .grid_clb_reset_E_out_out_2(resetWires[82]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[188]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[189]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[190]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[297]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[298]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[139]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[139]),
    .grid_clb_pReset_N_in_in_1(pResetWires[186]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[79]),
    .grid_clb_reset_W_in_in_1(resetWires[79]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[176]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[177]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[186]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[259]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[137]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[137]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__6_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_6_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_7__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__7_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__7_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__7_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__7_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[481]),
    .cby_config_enable_S_in_in_1(config_enableWires[481]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[282]),
    .grid_clb_pReset_N_in_in_2(pResetWires[533]),
    .grid_clb_Test_en_E_out_out_2(Test_enWires[236]),
    .grid_clb_reset_E_out_out_2(resetWires[236]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[202]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[203]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[533]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[318]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[319]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[159]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[159]),
    .grid_clb_pReset_N_in_in_1(pResetWires[529]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[233]),
    .grid_clb_reset_W_in_in_1(resetWires[233]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[162]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[163]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[529]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[280]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[157]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[157]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__7_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_7_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_9__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__8_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__8_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__8_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__8_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[146]),
    .cby_config_enable_S_in_in_1(config_enableWires[146]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[337]),
    .grid_clb_pReset_N_in_in_2(pResetWires[198]),
    .grid_clb_Test_en_E_out_out_2(Test_enWires[86]),
    .grid_clb_reset_E_out_out_2(resetWires[86]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[240]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[241]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[198]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[373]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[374]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[181]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[181]),
    .grid_clb_pReset_N_in_in_1(pResetWires[194]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[83]),
    .grid_clb_reset_W_in_in_1(resetWires[83]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[228]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[229]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[194]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[335]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[179]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[179]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__8_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_8_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_9__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__9_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__9_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__9_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__9_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[489]),
    .cby_config_enable_S_in_in_1(config_enableWires[489]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[358]),
    .grid_clb_pReset_N_in_in_2(pResetWires[541]),
    .grid_clb_Test_en_E_out_out_2(Test_enWires[240]),
    .grid_clb_reset_E_out_out_2(resetWires[240]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[254]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[255]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[541]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[394]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[395]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[201]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[201]),
    .grid_clb_pReset_N_in_in_1(pResetWires[537]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[237]),
    .grid_clb_reset_W_in_in_1(resetWires[237]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[214]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[215]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[537]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[356]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[199]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[199]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(cby_2__3__9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_9_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_11__3_
  (
    .cby_chany_top_out_out_1(cby_1__3__10_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__10_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__10_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__10_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[154]),
    .cby_config_enable_S_in_in_1(config_enableWires[154]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[413]),
    .grid_clb_pReset_N_in_in_2(pResetWires[206]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[292]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[293]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[206]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[449]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[450]),
    .grid_clb_prog_clk_0_N_in_in_2(prog_clk_1_wires[223]),
    .grid_clb_clk_0_N_in_in_2(clk_1_wires[223]),
    .grid_clb_pReset_N_in_in_1(pResetWires[202]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[87]),
    .grid_clb_reset_W_in_in_1(resetWires[87]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[280]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[281]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[202]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[411]),
    .grid_clb_prog_clk_0_N_in_in_1(prog_clk_1_wires[221]),
    .grid_clb_clk_0_N_in_in_1(clk_1_wires[221]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(grid_io_right_right_9_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_10_ccff_tail)
  );


  grid_mult_18
  grid_mult_18_11__10_
  (
    .cby_chany_top_out_out_1(cby_1__3__11_chany_top_out[0:19]),
    .cby_chany_bottom_out_out_1(cby_1__3__11_chany_bottom_out[0:19]),
    .cby_chany_top_in_in_1(sb_1__3__11_chany_bottom_out[0:19]),
    .cby_chany_bottom_in_in_1(sb_1__2__11_chany_top_out[0:19]),
    .cby_pReset_S_in_in_1(pResetWires[497]),
    .cby_config_enable_S_in_in_1(config_enableWires[497]),
    .cby_prog_clk_0_S_out_out_1(prog_clk_0_wires[434]),
    .grid_clb_pReset_N_in_in_2(pResetWires[549]),
    .grid_clb_sc_head_S_in_in_2(sc_headWires[306]),
    .grid_clb_sc_head_N_out_out_2(sc_headWires[307]),
    .grid_clb_config_enable_N_in_in_2(config_enableWires[549]),
    .grid_clb_prog_clk_0_S_out_out_2(prog_clk_0_wires[470]),
    .grid_clb_prog_clk_0_E_out_out_2(prog_clk_0_wires[471]),
    .grid_clb_prog_clk_0_S_in_in_2(prog_clk_1_wires[243]),
    .grid_clb_clk_0_S_in_in_2(clk_1_wires[243]),
    .grid_clb_pReset_N_in_in_1(pResetWires[545]),
    .grid_clb_Test_en_W_in_in_1(Test_enWires[241]),
    .grid_clb_reset_W_in_in_1(resetWires[241]),
    .grid_clb_sc_head_N_in_in_1(sc_headWires[266]),
    .grid_clb_sc_head_S_out_out_1(sc_headWires[267]),
    .grid_clb_config_enable_N_in_in_1(config_enableWires[545]),
    .grid_clb_prog_clk_0_S_out_out_1(prog_clk_0_wires[432]),
    .grid_clb_prog_clk_0_S_in_in_1(prog_clk_1_wires[241]),
    .grid_clb_clk_0_S_in_in_1(clk_1_wires[241]),
    .top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .right_width_1_height_0_subtile_0__pin_a_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .right_width_1_height_0_subtile_0__pin_a_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .right_width_1_height_0_subtile_0__pin_a_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .right_width_1_height_0_subtile_0__pin_a_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .right_width_1_height_0_subtile_0__pin_a_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .right_width_1_height_0_subtile_0__pin_a_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .right_width_1_height_0_subtile_0__pin_b_12_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .right_width_1_height_0_subtile_0__pin_b_13_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .right_width_1_height_0_subtile_0__pin_b_14_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .right_width_1_height_0_subtile_0__pin_b_15_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .right_width_1_height_0_subtile_0__pin_b_16_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .right_width_1_height_0_subtile_0__pin_b_17_(cby_12__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_head(grid_io_right_right_2_ccff_tail),
    .top_width_0_height_0_subtile_0__pin_out_0_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .top_width_0_height_0_subtile_0__pin_out_0_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .top_width_0_height_0_subtile_0__pin_out_1_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .top_width_0_height_0_subtile_0__pin_out_1_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .top_width_0_height_0_subtile_0__pin_out_2_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .top_width_0_height_0_subtile_0__pin_out_2_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .top_width_0_height_0_subtile_0__pin_out_3_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .top_width_0_height_0_subtile_0__pin_out_3_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .top_width_0_height_0_subtile_0__pin_out_4_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .top_width_0_height_0_subtile_0__pin_out_4_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .top_width_0_height_0_subtile_0__pin_out_5_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .top_width_0_height_0_subtile_0__pin_out_5_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .top_width_0_height_0_subtile_0__pin_out_6_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .top_width_0_height_0_subtile_0__pin_out_6_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .top_width_0_height_0_subtile_0__pin_out_7_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .top_width_0_height_0_subtile_0__pin_out_7_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .top_width_0_height_0_subtile_0__pin_out_8_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .top_width_0_height_0_subtile_0__pin_out_8_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .top_width_0_height_0_subtile_0__pin_out_9_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .top_width_0_height_0_subtile_0__pin_out_9_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .top_width_0_height_0_subtile_0__pin_out_10_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .top_width_0_height_0_subtile_0__pin_out_10_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .top_width_0_height_0_subtile_0__pin_out_11_upper(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .top_width_0_height_0_subtile_0__pin_out_11_lower(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .top_width_1_height_0_subtile_0__pin_out_12_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .top_width_1_height_0_subtile_0__pin_out_12_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .top_width_1_height_0_subtile_0__pin_out_13_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .top_width_1_height_0_subtile_0__pin_out_13_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .top_width_1_height_0_subtile_0__pin_out_14_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .top_width_1_height_0_subtile_0__pin_out_14_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .top_width_1_height_0_subtile_0__pin_out_15_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .top_width_1_height_0_subtile_0__pin_out_15_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .top_width_1_height_0_subtile_0__pin_out_16_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .top_width_1_height_0_subtile_0__pin_out_16_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .top_width_1_height_0_subtile_0__pin_out_17_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .top_width_1_height_0_subtile_0__pin_out_17_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .top_width_1_height_0_subtile_0__pin_out_18_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .top_width_1_height_0_subtile_0__pin_out_18_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .top_width_1_height_0_subtile_0__pin_out_19_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .top_width_1_height_0_subtile_0__pin_out_19_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .top_width_1_height_0_subtile_0__pin_out_20_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .top_width_1_height_0_subtile_0__pin_out_20_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .top_width_1_height_0_subtile_0__pin_out_21_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .top_width_1_height_0_subtile_0__pin_out_21_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .top_width_1_height_0_subtile_0__pin_out_22_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .top_width_1_height_0_subtile_0__pin_out_22_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .top_width_1_height_0_subtile_0__pin_out_23_upper(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .top_width_1_height_0_subtile_0__pin_out_23_lower(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .right_width_1_height_0_subtile_0__pin_out_24_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .right_width_1_height_0_subtile_0__pin_out_24_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .right_width_1_height_0_subtile_0__pin_out_25_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .right_width_1_height_0_subtile_0__pin_out_25_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .right_width_1_height_0_subtile_0__pin_out_26_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .right_width_1_height_0_subtile_0__pin_out_26_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .right_width_1_height_0_subtile_0__pin_out_27_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .right_width_1_height_0_subtile_0__pin_out_27_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .right_width_1_height_0_subtile_0__pin_out_28_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .right_width_1_height_0_subtile_0__pin_out_28_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .right_width_1_height_0_subtile_0__pin_out_29_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .right_width_1_height_0_subtile_0__pin_out_29_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .right_width_1_height_0_subtile_0__pin_out_30_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .right_width_1_height_0_subtile_0__pin_out_30_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .right_width_1_height_0_subtile_0__pin_out_31_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .right_width_1_height_0_subtile_0__pin_out_31_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .right_width_1_height_0_subtile_0__pin_out_32_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .right_width_1_height_0_subtile_0__pin_out_32_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .right_width_1_height_0_subtile_0__pin_out_33_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .right_width_1_height_0_subtile_0__pin_out_33_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .right_width_1_height_0_subtile_0__pin_out_34_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .right_width_1_height_0_subtile_0__pin_out_34_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .right_width_1_height_0_subtile_0__pin_out_35_upper(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .right_width_1_height_0_subtile_0__pin_out_35_lower(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .ccff_tail(grid_mult_18_11_ccff_tail)
  );


  sb_0__0_
  sb_0__0_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[5]),
    .config_enable_E_in(config_enableWires[25]),
    .pReset_E_in(pResetWires[25]),
    .chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_0_ccff_tail),
    .chany_top_out(sb_0__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
    .ccff_tail(sb_0__0__0_ccff_tail)
  );


  sb_0__1_
  sb_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[4]),
    .config_enable_S_out(config_enableWires[64]),
    .config_enable_E_in(config_enableWires[61]),
    .pReset_S_out(pResetWires[64]),
    .pReset_E_in(pResetWires[61]),
    .chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_1_ccff_tail),
    .chany_top_out(sb_0__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__0_ccff_tail)
  );


  sb_0__1_
  sb_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[10]),
    .config_enable_S_out(config_enableWires[113]),
    .config_enable_E_in(config_enableWires[110]),
    .pReset_S_out(pResetWires[113]),
    .pReset_E_in(pResetWires[110]),
    .chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_2_ccff_tail),
    .chany_top_out(sb_0__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__1_ccff_tail)
  );


  sb_0__1_
  sb_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[20]),
    .config_enable_S_out(config_enableWires[211]),
    .config_enable_E_in(config_enableWires[208]),
    .pReset_S_out(pResetWires[211]),
    .pReset_E_in(pResetWires[208]),
    .chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_4_ccff_tail),
    .chany_top_out(sb_0__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__2_ccff_tail)
  );


  sb_0__1_
  sb_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[25]),
    .config_enable_S_out(config_enableWires[260]),
    .config_enable_E_in(config_enableWires[257]),
    .pReset_S_out(pResetWires[260]),
    .pReset_E_in(pResetWires[257]),
    .chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_5_ccff_tail),
    .chany_top_out(sb_0__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__3_ccff_tail)
  );


  sb_0__1_
  sb_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[30]),
    .config_enable_S_out(config_enableWires[309]),
    .config_enable_E_in(config_enableWires[306]),
    .pReset_S_out(pResetWires[309]),
    .pReset_E_in(pResetWires[306]),
    .chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_6_ccff_tail),
    .chany_top_out(sb_0__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__4_ccff_tail)
  );


  sb_0__1_
  sb_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[35]),
    .config_enable_S_out(config_enableWires[358]),
    .config_enable_E_in(config_enableWires[355]),
    .pReset_S_out(pResetWires[358]),
    .pReset_E_in(pResetWires[355]),
    .chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_7_ccff_tail),
    .chany_top_out(sb_0__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__5_ccff_tail)
  );


  sb_0__1_
  sb_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[40]),
    .config_enable_S_out(config_enableWires[407]),
    .config_enable_E_in(config_enableWires[404]),
    .pReset_S_out(pResetWires[407]),
    .pReset_E_in(pResetWires[404]),
    .chany_top_in(cby_0__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_8_ccff_tail),
    .chany_top_out(sb_0__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__6_ccff_tail)
  );


  sb_0__1_
  sb_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[45]),
    .config_enable_S_out(config_enableWires[456]),
    .config_enable_E_in(config_enableWires[453]),
    .pReset_S_out(pResetWires[456]),
    .pReset_E_in(pResetWires[453]),
    .chany_top_in(cby_0__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_9_ccff_tail),
    .chany_top_out(sb_0__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__7_ccff_tail)
  );


  sb_0__1_
  sb_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[55]),
    .config_enable_S_out(config_enableWires[554]),
    .config_enable_E_in(config_enableWires[551]),
    .pReset_S_out(pResetWires[554]),
    .pReset_E_in(pResetWires[551]),
    .chany_top_in(cby_0__1__11_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__10_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_11_ccff_tail),
    .chany_top_out(sb_0__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__8_ccff_tail)
  );


  sb_0__3_
  sb_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[15]),
    .config_enable_S_out(config_enableWires[162]),
    .config_enable_E_in(config_enableWires[159]),
    .pReset_S_out(pResetWires[162]),
    .pReset_E_in(pResetWires[159]),
    .chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__3__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_3_ccff_tail),
    .chany_top_out(sb_0__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__3__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__3__0_ccff_tail)
  );


  sb_0__3_
  sb_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[50]),
    .config_enable_S_out(config_enableWires[505]),
    .config_enable_E_in(config_enableWires[502]),
    .pReset_S_out(pResetWires[505]),
    .pReset_E_in(pResetWires[502]),
    .chany_top_in(cby_0__1__10_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_right_in(cbx_1__3__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_0__1__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_left_left_10_ccff_tail),
    .chany_top_out(sb_0__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__3__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__3__1_ccff_tail)
  );


  sb_0__4_
  sb_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[62]),
    .config_enable_S_out(config_enableWires[603]),
    .config_enable_E_in(config_enableWires[600]),
    .sc_head_E_out(sc_headWires[1]),
    .sc_head_W_in(sc_head),
    .pReset_S_out(pResetWires[603]),
    .pReset_E_in(pResetWires[600]),
    .chanx_right_in(cbx_1__12__0_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_0__1__11_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .ccff_head(grid_io_top_top_0_ccff_tail),
    .chanx_right_out(sb_0__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__12__0_ccff_tail)
  );


  sb_1__0_
  sb_1__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[2]),
    .config_enable_E_in(config_enableWires[28]),
    .config_enable_N_out(config_enableWires[27]),
    .config_enable_W_out(config_enableWires[26]),
    .sc_head_E_out(sc_headWires[27]),
    .sc_head_W_in(sc_headWires[26]),
    .pReset_E_in(pResetWires[28]),
    .pReset_N_out(pResetWires[27]),
    .pReset_W_out(pResetWires[26]),
    .chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_11_ccff_tail),
    .chany_top_out(sb_1__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__0_ccff_tail)
  );


  sb_1__0_
  sb_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[65]),
    .config_enable_E_in(config_enableWires[31]),
    .config_enable_N_out(config_enableWires[30]),
    .config_enable_W_out(config_enableWires[29]),
    .pReset_E_in(pResetWires[31]),
    .pReset_N_out(pResetWires[30]),
    .pReset_W_out(pResetWires[29]),
    .chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_10_ccff_tail),
    .chany_top_out(sb_1__0__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__1_ccff_tail)
  );


  sb_1__0_
  sb_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[103]),
    .config_enable_E_in(config_enableWires[34]),
    .config_enable_N_out(config_enableWires[33]),
    .config_enable_W_out(config_enableWires[32]),
    .sc_head_E_out(sc_headWires[79]),
    .sc_head_W_in(sc_headWires[78]),
    .pReset_E_in(pResetWires[34]),
    .pReset_N_out(pResetWires[33]),
    .pReset_W_out(pResetWires[32]),
    .chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_9_ccff_tail),
    .chany_top_out(sb_1__0__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__2_ccff_tail)
  );


  sb_1__0_
  sb_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[141]),
    .config_enable_E_in(config_enableWires[37]),
    .config_enable_N_out(config_enableWires[36]),
    .config_enable_W_out(config_enableWires[35]),
    .pReset_E_in(pResetWires[37]),
    .pReset_N_out(pResetWires[36]),
    .pReset_W_out(pResetWires[35]),
    .chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_8_ccff_tail),
    .chany_top_out(sb_1__0__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__3_ccff_tail)
  );


  sb_1__0_
  sb_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[179]),
    .config_enable_E_in(config_enableWires[40]),
    .config_enable_N_out(config_enableWires[39]),
    .config_enable_W_out(config_enableWires[38]),
    .sc_head_E_out(sc_headWires[131]),
    .sc_head_W_in(sc_headWires[130]),
    .pReset_E_in(pResetWires[40]),
    .pReset_N_out(pResetWires[39]),
    .pReset_W_out(pResetWires[38]),
    .chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_7_ccff_tail),
    .chany_top_out(sb_1__0__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__4_ccff_tail)
  );


  sb_1__0_
  sb_6__0_
  (
    .clk_3_N_out(clk_3_wires[90]),
    .clk_3_S_in(clk0),
    .prog_clk_3_N_out(prog_clk_3_wires[90]),
    .prog_clk_3_S_in(prog_clk),
    .prog_clk_0_N_in(prog_clk_0_wires[217]),
    .config_enable_E_out(config_enableWires[43]),
    .config_enable_W_out(config_enableWires[41]),
    .config_enable_N_out(config_enableWires[42]),
    .config_enable_S_in(config_enable),
    .reset_N_out(resetWires[1]),
    .reset_S_in(reset),
    .Test_en_N_out(Test_enWires[1]),
    .Test_en_S_in(Test_en),
    .pReset_E_out(pResetWires[43]),
    .pReset_W_out(pResetWires[41]),
    .pReset_N_out(pResetWires[42]),
    .pReset_S_in(pReset),
    .chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_6_ccff_tail),
    .chany_top_out(sb_1__0__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__5_ccff_tail)
  );


  sb_1__0_
  sb_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[255]),
    .config_enable_E_out(config_enableWires[46]),
    .config_enable_N_out(config_enableWires[45]),
    .config_enable_W_in(config_enableWires[44]),
    .sc_head_E_out(sc_headWires[183]),
    .sc_head_W_in(sc_headWires[182]),
    .pReset_E_out(pResetWires[46]),
    .pReset_N_out(pResetWires[45]),
    .pReset_W_in(pResetWires[44]),
    .chany_top_in(cby_1__1__60_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_5_ccff_tail),
    .chany_top_out(sb_1__0__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__6_ccff_tail)
  );


  sb_1__0_
  sb_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[293]),
    .config_enable_E_out(config_enableWires[49]),
    .config_enable_N_out(config_enableWires[48]),
    .config_enable_W_in(config_enableWires[47]),
    .pReset_E_out(pResetWires[49]),
    .pReset_N_out(pResetWires[48]),
    .pReset_W_in(pResetWires[47]),
    .chany_top_in(cby_1__1__70_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_4_ccff_tail),
    .chany_top_out(sb_1__0__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__7_ccff_tail)
  );


  sb_1__0_
  sb_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[331]),
    .config_enable_E_out(config_enableWires[52]),
    .config_enable_N_out(config_enableWires[51]),
    .config_enable_W_in(config_enableWires[50]),
    .sc_head_E_out(sc_headWires[235]),
    .sc_head_W_in(sc_headWires[234]),
    .pReset_E_out(pResetWires[52]),
    .pReset_N_out(pResetWires[51]),
    .pReset_W_in(pResetWires[50]),
    .chany_top_in(cby_1__1__80_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_3_ccff_tail),
    .chany_top_out(sb_1__0__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__8_ccff_tail)
  );


  sb_1__0_
  sb_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[369]),
    .config_enable_E_out(config_enableWires[55]),
    .config_enable_N_out(config_enableWires[54]),
    .config_enable_W_in(config_enableWires[53]),
    .pReset_E_out(pResetWires[55]),
    .pReset_N_out(pResetWires[54]),
    .pReset_W_in(pResetWires[53]),
    .chany_top_in(cby_1__1__90_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_2_ccff_tail),
    .chany_top_out(sb_1__0__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__9_ccff_tail)
  );


  sb_1__0_
  sb_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[407]),
    .config_enable_E_out(config_enableWires[58]),
    .config_enable_N_out(config_enableWires[57]),
    .config_enable_W_in(config_enableWires[56]),
    .sc_head_E_out(sc_headWires[287]),
    .sc_head_W_in(sc_headWires[286]),
    .pReset_E_out(pResetWires[58]),
    .pReset_N_out(pResetWires[57]),
    .pReset_W_in(pResetWires[56]),
    .chany_top_in(cby_1__1__100_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__0__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .chanx_left_in(cbx_1__0__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_1_ccff_tail),
    .chany_top_out(sb_1__0__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__10_ccff_tail)
  );


  sb_1__1_
  sb_1__1_
  (
    .clk_1_N_in(clk_2_wires[4]),
    .clk_1_W_out(clk_1_wires[2]),
    .clk_1_E_out(clk_1_wires[1]),
    .prog_clk_1_N_in(prog_clk_2_wires[4]),
    .prog_clk_1_W_out(prog_clk_1_wires[2]),
    .prog_clk_1_E_out(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[8]),
    .config_enable_E_in(config_enableWires[66]),
    .config_enable_N_out(config_enableWires[65]),
    .config_enable_W_out(config_enableWires[62]),
    .pReset_E_in(pResetWires[66]),
    .pReset_N_out(pResetWires[65]),
    .pReset_W_out(pResetWires[62]),
    .chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__0_ccff_tail),
    .chany_top_out(sb_1__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__0_ccff_tail)
  );


  sb_1__1_
  sb_1__4_
  (
    .clk_2_S_out(clk_2_wires[10]),
    .clk_2_N_out(clk_2_wires[8]),
    .clk_2_E_in(clk_2_wires[6]),
    .prog_clk_2_S_out(prog_clk_2_wires[10]),
    .prog_clk_2_N_out(prog_clk_2_wires[8]),
    .prog_clk_2_E_in(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[23]),
    .config_enable_E_in(config_enableWires[213]),
    .config_enable_N_out(config_enableWires[212]),
    .config_enable_W_out(config_enableWires[209]),
    .pReset_E_in(pResetWires[213]),
    .pReset_N_out(pResetWires[212]),
    .pReset_W_out(pResetWires[209]),
    .chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__2_ccff_tail),
    .chany_top_out(sb_1__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__1_ccff_tail)
  );


  sb_1__1_
  sb_1__5_
  (
    .clk_1_S_in(clk_2_wires[9]),
    .clk_1_W_out(clk_1_wires[16]),
    .clk_1_E_out(clk_1_wires[15]),
    .prog_clk_1_S_in(prog_clk_2_wires[9]),
    .prog_clk_1_W_out(prog_clk_1_wires[16]),
    .prog_clk_1_E_out(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[28]),
    .config_enable_E_in(config_enableWires[262]),
    .config_enable_N_out(config_enableWires[261]),
    .config_enable_W_out(config_enableWires[258]),
    .pReset_E_in(pResetWires[262]),
    .pReset_N_out(pResetWires[261]),
    .pReset_W_out(pResetWires[258]),
    .chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__3_ccff_tail),
    .chany_top_out(sb_1__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__2_ccff_tail)
  );


  sb_1__1_
  sb_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[33]),
    .config_enable_E_in(config_enableWires[311]),
    .config_enable_N_out(config_enableWires[310]),
    .config_enable_W_out(config_enableWires[307]),
    .pReset_E_in(pResetWires[311]),
    .pReset_N_out(pResetWires[310]),
    .pReset_W_out(pResetWires[307]),
    .chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__4_ccff_tail),
    .chany_top_out(sb_1__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__3_ccff_tail)
  );


  sb_1__1_
  sb_1__7_
  (
    .clk_1_N_in(clk_2_wires[18]),
    .clk_1_W_out(clk_1_wires[23]),
    .clk_1_E_out(clk_1_wires[22]),
    .prog_clk_1_N_in(prog_clk_2_wires[18]),
    .prog_clk_1_W_out(prog_clk_1_wires[23]),
    .prog_clk_1_E_out(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[38]),
    .config_enable_E_in(config_enableWires[360]),
    .config_enable_N_out(config_enableWires[359]),
    .config_enable_W_out(config_enableWires[356]),
    .pReset_E_in(pResetWires[360]),
    .pReset_N_out(pResetWires[359]),
    .pReset_W_out(pResetWires[356]),
    .chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__5_ccff_tail),
    .chany_top_out(sb_1__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__4_ccff_tail)
  );


  sb_1__1_
  sb_1__8_
  (
    .clk_2_S_out(clk_2_wires[17]),
    .clk_2_N_out(clk_2_wires[15]),
    .clk_2_E_in(clk_2_wires[13]),
    .prog_clk_2_S_out(prog_clk_2_wires[17]),
    .prog_clk_2_N_out(prog_clk_2_wires[15]),
    .prog_clk_2_E_in(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[43]),
    .config_enable_E_in(config_enableWires[409]),
    .config_enable_N_out(config_enableWires[408]),
    .config_enable_W_out(config_enableWires[405]),
    .pReset_E_in(pResetWires[409]),
    .pReset_N_out(pResetWires[408]),
    .pReset_W_out(pResetWires[405]),
    .chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__6_ccff_tail),
    .chany_top_out(sb_1__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__5_ccff_tail)
  );


  sb_1__1_
  sb_1__11_
  (
    .clk_1_S_in(clk_2_wires[23]),
    .clk_1_W_out(clk_1_wires[37]),
    .clk_1_E_out(clk_1_wires[36]),
    .prog_clk_1_S_in(prog_clk_2_wires[23]),
    .prog_clk_1_W_out(prog_clk_1_wires[37]),
    .prog_clk_1_E_out(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[58]),
    .config_enable_E_in(config_enableWires[556]),
    .config_enable_N_out(config_enableWires[555]),
    .config_enable_W_out(config_enableWires[552]),
    .pReset_E_in(pResetWires[556]),
    .pReset_N_out(pResetWires[555]),
    .pReset_W_out(pResetWires[552]),
    .chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__8_ccff_tail),
    .chany_top_out(sb_1__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__6_ccff_tail)
  );


  sb_1__1_
  sb_2__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[68]),
    .config_enable_E_in(config_enableWires[70]),
    .config_enable_N_out(config_enableWires[69]),
    .config_enable_W_out(config_enableWires[67]),
    .pReset_E_in(pResetWires[70]),
    .pReset_N_out(pResetWires[69]),
    .pReset_W_out(pResetWires[67]),
    .chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__9_ccff_tail),
    .chany_top_out(sb_1__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__7_ccff_tail)
  );


  sb_1__1_
  sb_2__4_
  (
    .clk_3_S_out(clk_3_wires[64]),
    .clk_2_N_in(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[59]),
    .clk_2_W_out(clk_2_wires[7]),
    .prog_clk_3_S_out(prog_clk_3_wires[64]),
    .prog_clk_2_N_in(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[59]),
    .prog_clk_2_W_out(prog_clk_2_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[77]),
    .config_enable_E_in(config_enableWires[217]),
    .config_enable_N_out(config_enableWires[216]),
    .config_enable_W_out(config_enableWires[214]),
    .pReset_E_in(pResetWires[217]),
    .pReset_N_out(pResetWires[216]),
    .pReset_W_out(pResetWires[214]),
    .chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__11_ccff_tail),
    .chany_top_out(sb_1__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__8_ccff_tail)
  );


  sb_1__1_
  sb_2__5_
  (
    .clk_3_S_out(clk_3_wires[58]),
    .clk_3_N_in(clk_3_wires[55]),
    .prog_clk_3_S_out(prog_clk_3_wires[58]),
    .prog_clk_3_N_in(prog_clk_3_wires[55]),
    .prog_clk_0_N_in(prog_clk_0_wires[80]),
    .config_enable_E_in(config_enableWires[266]),
    .config_enable_N_out(config_enableWires[265]),
    .config_enable_W_out(config_enableWires[263]),
    .pReset_E_in(pResetWires[266]),
    .pReset_N_out(pResetWires[265]),
    .pReset_W_out(pResetWires[263]),
    .chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__12_ccff_tail),
    .chany_top_out(sb_1__1__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__9_ccff_tail)
  );


  sb_1__1_
  sb_2__6_
  (
    .clk_3_S_out(clk_3_wires[54]),
    .clk_3_N_out(clk_3_wires[52]),
    .clk_3_E_in(clk_3_wires[51]),
    .prog_clk_3_S_out(prog_clk_3_wires[54]),
    .prog_clk_3_N_out(prog_clk_3_wires[52]),
    .prog_clk_3_E_in(prog_clk_3_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[83]),
    .config_enable_E_in(config_enableWires[315]),
    .config_enable_N_out(config_enableWires[314]),
    .config_enable_W_out(config_enableWires[312]),
    .pReset_E_in(pResetWires[315]),
    .pReset_N_out(pResetWires[314]),
    .pReset_W_out(pResetWires[312]),
    .chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__13_ccff_tail),
    .chany_top_out(sb_1__1__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__10_ccff_tail)
  );


  sb_1__1_
  sb_2__7_
  (
    .clk_3_N_out(clk_3_wires[56]),
    .clk_3_S_in(clk_3_wires[53]),
    .prog_clk_3_N_out(prog_clk_3_wires[56]),
    .prog_clk_3_S_in(prog_clk_3_wires[53]),
    .prog_clk_0_N_in(prog_clk_0_wires[86]),
    .config_enable_E_in(config_enableWires[364]),
    .config_enable_N_out(config_enableWires[363]),
    .config_enable_W_out(config_enableWires[361]),
    .pReset_E_in(pResetWires[364]),
    .pReset_N_out(pResetWires[363]),
    .pReset_W_out(pResetWires[361]),
    .chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__14_ccff_tail),
    .chany_top_out(sb_1__1__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__11_ccff_tail)
  );


  sb_1__1_
  sb_2__8_
  (
    .clk_3_N_out(clk_3_wires[62]),
    .clk_2_S_in(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[57]),
    .clk_2_W_out(clk_2_wires[14]),
    .prog_clk_3_N_out(prog_clk_3_wires[62]),
    .prog_clk_2_S_in(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[57]),
    .prog_clk_2_W_out(prog_clk_2_wires[14]),
    .prog_clk_0_N_in(prog_clk_0_wires[89]),
    .config_enable_E_in(config_enableWires[413]),
    .config_enable_N_out(config_enableWires[412]),
    .config_enable_W_out(config_enableWires[410]),
    .pReset_E_in(pResetWires[413]),
    .pReset_N_out(pResetWires[412]),
    .pReset_W_out(pResetWires[410]),
    .chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__15_ccff_tail),
    .chany_top_out(sb_1__1__12_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__12_ccff_tail)
  );


  sb_1__1_
  sb_2__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[98]),
    .config_enable_E_in(config_enableWires[560]),
    .config_enable_N_out(config_enableWires[559]),
    .config_enable_W_out(config_enableWires[557]),
    .pReset_E_in(pResetWires[560]),
    .pReset_N_out(pResetWires[559]),
    .pReset_W_out(pResetWires[557]),
    .chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__17_ccff_tail),
    .chany_top_out(sb_1__1__13_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__13_ccff_tail)
  );


  sb_1__1_
  sb_3__1_
  (
    .clk_1_N_in(clk_2_wires[30]),
    .clk_1_W_out(clk_1_wires[44]),
    .clk_1_E_out(clk_1_wires[43]),
    .prog_clk_1_N_in(prog_clk_2_wires[30]),
    .prog_clk_1_W_out(prog_clk_1_wires[44]),
    .prog_clk_1_E_out(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[106]),
    .config_enable_E_in(config_enableWires[74]),
    .config_enable_N_out(config_enableWires[73]),
    .config_enable_W_out(config_enableWires[71]),
    .pReset_E_in(pResetWires[74]),
    .pReset_N_out(pResetWires[73]),
    .pReset_W_out(pResetWires[71]),
    .chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__18_ccff_tail),
    .chany_top_out(sb_1__1__14_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__14_ccff_tail)
  );


  sb_1__1_
  sb_3__4_
  (
    .clk_2_S_out(clk_2_wires[40]),
    .clk_2_N_out(clk_2_wires[38]),
    .clk_2_E_in(clk_2_wires[37]),
    .prog_clk_2_S_out(prog_clk_2_wires[40]),
    .prog_clk_2_N_out(prog_clk_2_wires[38]),
    .prog_clk_2_E_in(prog_clk_2_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[115]),
    .config_enable_E_in(config_enableWires[221]),
    .config_enable_N_out(config_enableWires[220]),
    .config_enable_W_out(config_enableWires[218]),
    .pReset_E_in(pResetWires[221]),
    .pReset_N_out(pResetWires[220]),
    .pReset_W_out(pResetWires[218]),
    .chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__20_ccff_tail),
    .chany_top_out(sb_1__1__15_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__15_ccff_tail)
  );


  sb_1__1_
  sb_3__5_
  (
    .clk_1_S_in(clk_2_wires[39]),
    .clk_1_W_out(clk_1_wires[58]),
    .clk_1_E_out(clk_1_wires[57]),
    .prog_clk_1_S_in(prog_clk_2_wires[39]),
    .prog_clk_1_W_out(prog_clk_1_wires[58]),
    .prog_clk_1_E_out(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[118]),
    .config_enable_E_in(config_enableWires[270]),
    .config_enable_N_out(config_enableWires[269]),
    .config_enable_W_out(config_enableWires[267]),
    .pReset_E_in(pResetWires[270]),
    .pReset_N_out(pResetWires[269]),
    .pReset_W_out(pResetWires[267]),
    .chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__21_ccff_tail),
    .chany_top_out(sb_1__1__16_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__16_ccff_tail)
  );


  sb_1__1_
  sb_3__6_
  (
    .clk_3_W_out(clk_3_wires[50]),
    .clk_3_E_in(clk_3_wires[47]),
    .prog_clk_3_W_out(prog_clk_3_wires[50]),
    .prog_clk_3_E_in(prog_clk_3_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[121]),
    .config_enable_E_in(config_enableWires[319]),
    .config_enable_N_out(config_enableWires[318]),
    .config_enable_W_out(config_enableWires[316]),
    .pReset_E_in(pResetWires[319]),
    .pReset_N_out(pResetWires[318]),
    .pReset_W_out(pResetWires[316]),
    .chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__22_ccff_tail),
    .chany_top_out(sb_1__1__17_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__17_ccff_tail)
  );


  sb_1__1_
  sb_3__7_
  (
    .clk_1_N_in(clk_2_wires[54]),
    .clk_1_W_out(clk_1_wires[65]),
    .clk_1_E_out(clk_1_wires[64]),
    .prog_clk_1_N_in(prog_clk_2_wires[54]),
    .prog_clk_1_W_out(prog_clk_1_wires[65]),
    .prog_clk_1_E_out(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[124]),
    .config_enable_E_in(config_enableWires[368]),
    .config_enable_N_out(config_enableWires[367]),
    .config_enable_W_out(config_enableWires[365]),
    .pReset_E_in(pResetWires[368]),
    .pReset_N_out(pResetWires[367]),
    .pReset_W_out(pResetWires[365]),
    .chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__23_ccff_tail),
    .chany_top_out(sb_1__1__18_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__18_ccff_tail)
  );


  sb_1__1_
  sb_3__8_
  (
    .clk_2_S_out(clk_2_wires[53]),
    .clk_2_N_out(clk_2_wires[51]),
    .clk_2_E_in(clk_2_wires[50]),
    .prog_clk_2_S_out(prog_clk_2_wires[53]),
    .prog_clk_2_N_out(prog_clk_2_wires[51]),
    .prog_clk_2_E_in(prog_clk_2_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[127]),
    .config_enable_E_in(config_enableWires[417]),
    .config_enable_N_out(config_enableWires[416]),
    .config_enable_W_out(config_enableWires[414]),
    .pReset_E_in(pResetWires[417]),
    .pReset_N_out(pResetWires[416]),
    .pReset_W_out(pResetWires[414]),
    .chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__24_ccff_tail),
    .chany_top_out(sb_1__1__19_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__19_ccff_tail)
  );


  sb_1__1_
  sb_3__11_
  (
    .clk_1_S_in(clk_2_wires[65]),
    .clk_1_W_out(clk_1_wires[79]),
    .clk_1_E_out(clk_1_wires[78]),
    .prog_clk_1_S_in(prog_clk_2_wires[65]),
    .prog_clk_1_W_out(prog_clk_1_wires[79]),
    .prog_clk_1_E_out(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[136]),
    .config_enable_E_in(config_enableWires[564]),
    .config_enable_N_out(config_enableWires[563]),
    .config_enable_W_out(config_enableWires[561]),
    .pReset_E_in(pResetWires[564]),
    .pReset_N_out(pResetWires[563]),
    .pReset_W_out(pResetWires[561]),
    .chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__26_ccff_tail),
    .chany_top_out(sb_1__1__20_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__20_ccff_tail)
  );


  sb_1__1_
  sb_4__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[144]),
    .config_enable_E_in(config_enableWires[78]),
    .config_enable_N_out(config_enableWires[77]),
    .config_enable_W_out(config_enableWires[75]),
    .pReset_E_in(pResetWires[78]),
    .pReset_N_out(pResetWires[77]),
    .pReset_W_out(pResetWires[75]),
    .chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__27_ccff_tail),
    .chany_top_out(sb_1__1__21_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__21_ccff_tail)
  );


  sb_1__1_
  sb_4__4_
  (
    .clk_3_S_out(clk_3_wires[20]),
    .clk_2_N_in(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[15]),
    .clk_2_W_out(clk_2_wires[36]),
    .clk_2_E_out(clk_2_wires[34]),
    .prog_clk_3_S_out(prog_clk_3_wires[20]),
    .prog_clk_2_N_in(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[15]),
    .prog_clk_2_W_out(prog_clk_2_wires[36]),
    .prog_clk_2_E_out(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[153]),
    .config_enable_E_in(config_enableWires[225]),
    .config_enable_N_out(config_enableWires[224]),
    .config_enable_W_out(config_enableWires[222]),
    .pReset_E_in(pResetWires[225]),
    .pReset_N_out(pResetWires[224]),
    .pReset_W_out(pResetWires[222]),
    .chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__29_ccff_tail),
    .chany_top_out(sb_1__1__22_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__22_ccff_tail)
  );


  sb_1__1_
  sb_4__5_
  (
    .clk_3_S_out(clk_3_wires[14]),
    .clk_3_N_in(clk_3_wires[11]),
    .prog_clk_3_S_out(prog_clk_3_wires[14]),
    .prog_clk_3_N_in(prog_clk_3_wires[11]),
    .prog_clk_0_N_in(prog_clk_0_wires[156]),
    .config_enable_E_in(config_enableWires[274]),
    .config_enable_N_out(config_enableWires[273]),
    .config_enable_W_out(config_enableWires[271]),
    .pReset_E_in(pResetWires[274]),
    .pReset_N_out(pResetWires[273]),
    .pReset_W_out(pResetWires[271]),
    .chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__30_ccff_tail),
    .chany_top_out(sb_1__1__23_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__23_ccff_tail)
  );


  sb_1__1_
  sb_4__6_
  (
    .clk_3_W_out(clk_3_wires[46]),
    .clk_3_S_out(clk_3_wires[10]),
    .clk_3_N_out(clk_3_wires[8]),
    .clk_3_E_in(clk_3_wires[7]),
    .prog_clk_3_W_out(prog_clk_3_wires[46]),
    .prog_clk_3_S_out(prog_clk_3_wires[10]),
    .prog_clk_3_N_out(prog_clk_3_wires[8]),
    .prog_clk_3_E_in(prog_clk_3_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[159]),
    .config_enable_E_in(config_enableWires[323]),
    .config_enable_N_out(config_enableWires[322]),
    .config_enable_W_out(config_enableWires[320]),
    .pReset_E_in(pResetWires[323]),
    .pReset_N_out(pResetWires[322]),
    .pReset_W_out(pResetWires[320]),
    .chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__31_ccff_tail),
    .chany_top_out(sb_1__1__24_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__24_ccff_tail)
  );


  sb_1__1_
  sb_4__7_
  (
    .clk_3_N_out(clk_3_wires[12]),
    .clk_3_S_in(clk_3_wires[9]),
    .prog_clk_3_N_out(prog_clk_3_wires[12]),
    .prog_clk_3_S_in(prog_clk_3_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[162]),
    .config_enable_E_in(config_enableWires[372]),
    .config_enable_N_out(config_enableWires[371]),
    .config_enable_W_out(config_enableWires[369]),
    .pReset_E_in(pResetWires[372]),
    .pReset_N_out(pResetWires[371]),
    .pReset_W_out(pResetWires[369]),
    .chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__32_ccff_tail),
    .chany_top_out(sb_1__1__25_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__25_ccff_tail)
  );


  sb_1__1_
  sb_4__8_
  (
    .clk_3_N_out(clk_3_wires[18]),
    .clk_2_S_in(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[13]),
    .clk_2_W_out(clk_2_wires[49]),
    .clk_2_E_out(clk_2_wires[47]),
    .prog_clk_3_N_out(prog_clk_3_wires[18]),
    .prog_clk_2_S_in(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[13]),
    .prog_clk_2_W_out(prog_clk_2_wires[49]),
    .prog_clk_2_E_out(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[165]),
    .config_enable_E_in(config_enableWires[421]),
    .config_enable_N_out(config_enableWires[420]),
    .config_enable_W_out(config_enableWires[418]),
    .pReset_E_in(pResetWires[421]),
    .pReset_N_out(pResetWires[420]),
    .pReset_W_out(pResetWires[418]),
    .chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__33_ccff_tail),
    .chany_top_out(sb_1__1__26_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__26_ccff_tail)
  );


  sb_1__1_
  sb_4__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[174]),
    .config_enable_E_in(config_enableWires[568]),
    .config_enable_N_out(config_enableWires[567]),
    .config_enable_W_out(config_enableWires[565]),
    .pReset_E_in(pResetWires[568]),
    .pReset_N_out(pResetWires[567]),
    .pReset_W_out(pResetWires[565]),
    .chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__35_ccff_tail),
    .chany_top_out(sb_1__1__27_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__27_ccff_tail)
  );


  sb_1__1_
  sb_5__1_
  (
    .clk_1_N_in(clk_2_wires[32]),
    .clk_1_W_out(clk_1_wires[86]),
    .clk_1_E_out(clk_1_wires[85]),
    .prog_clk_1_N_in(prog_clk_2_wires[32]),
    .prog_clk_1_W_out(prog_clk_1_wires[86]),
    .prog_clk_1_E_out(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[182]),
    .config_enable_E_in(config_enableWires[82]),
    .config_enable_N_out(config_enableWires[81]),
    .config_enable_W_out(config_enableWires[79]),
    .pReset_E_in(pResetWires[82]),
    .pReset_N_out(pResetWires[81]),
    .pReset_W_out(pResetWires[79]),
    .chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__36_ccff_tail),
    .chany_top_out(sb_1__1__28_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__28_ccff_tail)
  );


  sb_1__1_
  sb_5__4_
  (
    .clk_2_S_out(clk_2_wires[44]),
    .clk_2_N_out(clk_2_wires[42]),
    .clk_2_W_in(clk_2_wires[35]),
    .prog_clk_2_S_out(prog_clk_2_wires[44]),
    .prog_clk_2_N_out(prog_clk_2_wires[42]),
    .prog_clk_2_W_in(prog_clk_2_wires[35]),
    .prog_clk_0_N_in(prog_clk_0_wires[191]),
    .config_enable_E_in(config_enableWires[229]),
    .config_enable_N_out(config_enableWires[228]),
    .config_enable_W_out(config_enableWires[226]),
    .pReset_E_in(pResetWires[229]),
    .pReset_N_out(pResetWires[228]),
    .pReset_W_out(pResetWires[226]),
    .chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__38_ccff_tail),
    .chany_top_out(sb_1__1__29_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__29_ccff_tail)
  );


  sb_1__1_
  sb_5__5_
  (
    .clk_1_S_in(clk_2_wires[43]),
    .clk_1_W_out(clk_1_wires[100]),
    .clk_1_E_out(clk_1_wires[99]),
    .prog_clk_1_S_in(prog_clk_2_wires[43]),
    .prog_clk_1_W_out(prog_clk_1_wires[100]),
    .prog_clk_1_E_out(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[194]),
    .config_enable_E_in(config_enableWires[278]),
    .config_enable_N_out(config_enableWires[277]),
    .config_enable_W_out(config_enableWires[275]),
    .pReset_E_in(pResetWires[278]),
    .pReset_N_out(pResetWires[277]),
    .pReset_W_out(pResetWires[275]),
    .chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__39_ccff_tail),
    .chany_top_out(sb_1__1__30_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__30_ccff_tail)
  );


  sb_1__1_
  sb_5__6_
  (
    .clk_3_W_out(clk_3_wires[6]),
    .clk_3_E_in(clk_3_wires[3]),
    .prog_clk_3_W_out(prog_clk_3_wires[6]),
    .prog_clk_3_E_in(prog_clk_3_wires[3]),
    .prog_clk_0_N_in(prog_clk_0_wires[197]),
    .config_enable_E_in(config_enableWires[327]),
    .config_enable_N_out(config_enableWires[326]),
    .config_enable_W_out(config_enableWires[324]),
    .pReset_E_in(pResetWires[327]),
    .pReset_N_out(pResetWires[326]),
    .pReset_W_out(pResetWires[324]),
    .chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__40_ccff_tail),
    .chany_top_out(sb_1__1__31_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__31_ccff_tail)
  );


  sb_1__1_
  sb_5__7_
  (
    .clk_1_N_in(clk_2_wires[58]),
    .clk_1_W_out(clk_1_wires[107]),
    .clk_1_E_out(clk_1_wires[106]),
    .prog_clk_1_N_in(prog_clk_2_wires[58]),
    .prog_clk_1_W_out(prog_clk_1_wires[107]),
    .prog_clk_1_E_out(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[200]),
    .config_enable_E_in(config_enableWires[376]),
    .config_enable_N_out(config_enableWires[375]),
    .config_enable_W_out(config_enableWires[373]),
    .pReset_E_in(pResetWires[376]),
    .pReset_N_out(pResetWires[375]),
    .pReset_W_out(pResetWires[373]),
    .chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__41_ccff_tail),
    .chany_top_out(sb_1__1__32_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__32_ccff_tail)
  );


  sb_1__1_
  sb_5__8_
  (
    .clk_2_S_out(clk_2_wires[57]),
    .clk_2_N_out(clk_2_wires[55]),
    .clk_2_W_in(clk_2_wires[48]),
    .prog_clk_2_S_out(prog_clk_2_wires[57]),
    .prog_clk_2_N_out(prog_clk_2_wires[55]),
    .prog_clk_2_W_in(prog_clk_2_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[203]),
    .config_enable_E_in(config_enableWires[425]),
    .config_enable_N_out(config_enableWires[424]),
    .config_enable_W_out(config_enableWires[422]),
    .pReset_E_in(pResetWires[425]),
    .pReset_N_out(pResetWires[424]),
    .pReset_W_out(pResetWires[422]),
    .chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__42_ccff_tail),
    .chany_top_out(sb_1__1__33_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__33_ccff_tail)
  );


  sb_1__1_
  sb_5__11_
  (
    .clk_1_S_in(clk_2_wires[67]),
    .clk_1_W_out(clk_1_wires[121]),
    .clk_1_E_out(clk_1_wires[120]),
    .prog_clk_1_S_in(prog_clk_2_wires[67]),
    .prog_clk_1_W_out(prog_clk_1_wires[121]),
    .prog_clk_1_E_out(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[212]),
    .config_enable_E_in(config_enableWires[572]),
    .config_enable_N_out(config_enableWires[571]),
    .config_enable_W_out(config_enableWires[569]),
    .pReset_E_in(pResetWires[572]),
    .pReset_N_out(pResetWires[571]),
    .pReset_W_out(pResetWires[569]),
    .chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__44_ccff_tail),
    .chany_top_out(sb_1__1__34_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__34_ccff_tail)
  );


  sb_1__1_
  sb_6__1_
  (
    .clk_3_N_out(clk_3_wires[92]),
    .clk_3_S_in(clk_3_wires[89]),
    .prog_clk_3_N_out(prog_clk_3_wires[92]),
    .prog_clk_3_S_in(prog_clk_3_wires[89]),
    .prog_clk_0_N_in(prog_clk_0_wires[220]),
    .config_enable_E_out(config_enableWires[86]),
    .config_enable_W_out(config_enableWires[83]),
    .config_enable_N_out(config_enableWires[85]),
    .config_enable_S_in(config_enableWires[2]),
    .reset_N_out(resetWires[3]),
    .reset_S_in(resetWires[2]),
    .Test_en_N_out(Test_enWires[3]),
    .Test_en_S_in(Test_enWires[2]),
    .pReset_E_out(pResetWires[86]),
    .pReset_W_out(pResetWires[83]),
    .pReset_N_out(pResetWires[85]),
    .pReset_S_in(pResetWires[2]),
    .chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__45_ccff_tail),
    .chany_top_out(sb_1__1__35_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__35_ccff_tail)
  );


  sb_1__1_
  sb_6__4_
  (
    .clk_3_N_out(clk_3_wires[98]),
    .clk_3_S_in(clk_3_wires[95]),
    .prog_clk_3_N_out(prog_clk_3_wires[98]),
    .prog_clk_3_S_in(prog_clk_3_wires[95]),
    .prog_clk_0_N_in(prog_clk_0_wires[229]),
    .config_enable_E_out(config_enableWires[233]),
    .config_enable_W_out(config_enableWires[230]),
    .config_enable_N_out(config_enableWires[232]),
    .config_enable_S_in(config_enableWires[8]),
    .reset_N_out(resetWires[9]),
    .reset_S_in(resetWires[8]),
    .Test_en_N_out(Test_enWires[9]),
    .Test_en_S_in(Test_enWires[8]),
    .pReset_E_out(pResetWires[233]),
    .pReset_W_out(pResetWires[230]),
    .pReset_N_out(pResetWires[232]),
    .pReset_S_in(pResetWires[8]),
    .chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__56_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__47_ccff_tail),
    .chany_top_out(sb_1__1__36_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__36_ccff_tail)
  );


  sb_1__1_
  sb_6__5_
  (
    .clk_3_N_out(clk_3_wires[100]),
    .clk_3_S_in(clk_3_wires[97]),
    .prog_clk_3_N_out(prog_clk_3_wires[100]),
    .prog_clk_3_S_in(prog_clk_3_wires[97]),
    .prog_clk_0_N_in(prog_clk_0_wires[232]),
    .config_enable_E_out(config_enableWires[282]),
    .config_enable_W_out(config_enableWires[279]),
    .config_enable_N_out(config_enableWires[281]),
    .config_enable_S_in(config_enableWires[10]),
    .reset_N_out(resetWires[11]),
    .reset_S_in(resetWires[10]),
    .Test_en_N_out(Test_enWires[11]),
    .Test_en_S_in(Test_enWires[10]),
    .pReset_E_out(pResetWires[282]),
    .pReset_W_out(pResetWires[279]),
    .pReset_N_out(pResetWires[281]),
    .pReset_S_in(pResetWires[10]),
    .chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__57_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__48_ccff_tail),
    .chany_top_out(sb_1__1__37_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__37_ccff_tail)
  );


  sb_1__1_
  sb_6__6_
  (
    .clk_3_S_in(clk_3_wires[99]),
    .clk_3_W_out(clk_3_wires[2]),
    .clk_3_E_out(clk_3_wires[0]),
    .prog_clk_3_S_in(prog_clk_3_wires[99]),
    .prog_clk_3_W_out(prog_clk_3_wires[2]),
    .prog_clk_3_E_out(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[235]),
    .config_enable_E_out(config_enableWires[331]),
    .config_enable_W_out(config_enableWires[328]),
    .config_enable_N_out(config_enableWires[330]),
    .config_enable_S_in(config_enableWires[12]),
    .reset_N_out(resetWires[13]),
    .reset_S_in(resetWires[12]),
    .Test_en_N_out(Test_enWires[13]),
    .Test_en_S_in(Test_enWires[12]),
    .pReset_E_out(pResetWires[331]),
    .pReset_W_out(pResetWires[328]),
    .pReset_N_out(pResetWires[330]),
    .pReset_S_in(pResetWires[12]),
    .chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__58_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__49_ccff_tail),
    .chany_top_out(sb_1__1__38_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__38_ccff_tail)
  );


  sb_1__1_
  sb_6__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[238]),
    .config_enable_E_out(config_enableWires[380]),
    .config_enable_W_out(config_enableWires[377]),
    .config_enable_N_out(config_enableWires[379]),
    .config_enable_S_in(config_enableWires[14]),
    .reset_N_out(resetWires[15]),
    .reset_S_in(resetWires[14]),
    .Test_en_N_out(Test_enWires[15]),
    .Test_en_S_in(Test_enWires[14]),
    .pReset_E_out(pResetWires[380]),
    .pReset_W_out(pResetWires[377]),
    .pReset_N_out(pResetWires[379]),
    .pReset_S_in(pResetWires[14]),
    .chany_top_in(cby_1__1__56_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__59_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__50_ccff_tail),
    .chany_top_out(sb_1__1__39_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__39_ccff_tail)
  );


  sb_1__1_
  sb_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[241]),
    .config_enable_E_out(config_enableWires[429]),
    .config_enable_W_out(config_enableWires[426]),
    .config_enable_N_out(config_enableWires[428]),
    .config_enable_S_in(config_enableWires[16]),
    .reset_N_out(resetWires[17]),
    .reset_S_in(resetWires[16]),
    .Test_en_N_out(Test_enWires[17]),
    .Test_en_S_in(Test_enWires[16]),
    .pReset_E_out(pResetWires[429]),
    .pReset_W_out(pResetWires[426]),
    .pReset_N_out(pResetWires[428]),
    .pReset_S_in(pResetWires[16]),
    .chany_top_in(cby_1__1__57_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__60_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__56_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__51_ccff_tail),
    .chany_top_out(sb_1__1__40_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__40_ccff_tail)
  );


  sb_1__1_
  sb_6__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[250]),
    .config_enable_E_out(config_enableWires[576]),
    .config_enable_W_out(config_enableWires[573]),
    .config_enable_N_out(config_enableWires[575]),
    .config_enable_S_in(config_enableWires[22]),
    .reset_N_out(resetWires[23]),
    .reset_S_in(resetWires[22]),
    .Test_en_N_out(Test_enWires[23]),
    .Test_en_S_in(Test_enWires[22]),
    .pReset_E_out(pResetWires[576]),
    .pReset_W_out(pResetWires[573]),
    .pReset_N_out(pResetWires[575]),
    .pReset_S_in(pResetWires[22]),
    .chany_top_in(cby_1__1__59_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__62_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__58_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__53_ccff_tail),
    .chany_top_out(sb_1__1__41_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__41_ccff_tail)
  );


  sb_1__1_
  sb_7__1_
  (
    .clk_1_N_in(clk_2_wires[74]),
    .clk_1_W_out(clk_1_wires[128]),
    .clk_1_E_out(clk_1_wires[127]),
    .prog_clk_1_N_in(prog_clk_2_wires[74]),
    .prog_clk_1_W_out(prog_clk_1_wires[128]),
    .prog_clk_1_E_out(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[258]),
    .config_enable_E_out(config_enableWires[90]),
    .config_enable_N_out(config_enableWires[89]),
    .config_enable_W_in(config_enableWires[87]),
    .pReset_E_out(pResetWires[90]),
    .pReset_N_out(pResetWires[89]),
    .pReset_W_in(pResetWires[87]),
    .chany_top_in(cby_1__1__61_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__63_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__60_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__54_ccff_tail),
    .chany_top_out(sb_1__1__42_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__42_ccff_tail)
  );


  sb_1__1_
  sb_7__4_
  (
    .clk_2_S_out(clk_2_wires[84]),
    .clk_2_N_out(clk_2_wires[82]),
    .clk_2_E_in(clk_2_wires[81]),
    .prog_clk_2_S_out(prog_clk_2_wires[84]),
    .prog_clk_2_N_out(prog_clk_2_wires[82]),
    .prog_clk_2_E_in(prog_clk_2_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[267]),
    .config_enable_E_out(config_enableWires[237]),
    .config_enable_N_out(config_enableWires[236]),
    .config_enable_W_in(config_enableWires[234]),
    .pReset_E_out(pResetWires[237]),
    .pReset_N_out(pResetWires[236]),
    .pReset_W_in(pResetWires[234]),
    .chany_top_in(cby_1__1__63_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__65_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__62_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__56_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__56_ccff_tail),
    .chany_top_out(sb_1__1__43_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__43_ccff_tail)
  );


  sb_1__1_
  sb_7__5_
  (
    .clk_1_S_in(clk_2_wires[83]),
    .clk_1_W_out(clk_1_wires[142]),
    .clk_1_E_out(clk_1_wires[141]),
    .prog_clk_1_S_in(prog_clk_2_wires[83]),
    .prog_clk_1_W_out(prog_clk_1_wires[142]),
    .prog_clk_1_E_out(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[270]),
    .config_enable_E_out(config_enableWires[286]),
    .config_enable_N_out(config_enableWires[285]),
    .config_enable_W_in(config_enableWires[283]),
    .pReset_E_out(pResetWires[286]),
    .pReset_N_out(pResetWires[285]),
    .pReset_W_in(pResetWires[283]),
    .chany_top_in(cby_1__1__64_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__66_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__63_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__57_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__57_ccff_tail),
    .chany_top_out(sb_1__1__44_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__44_ccff_tail)
  );


  sb_1__1_
  sb_7__6_
  (
    .clk_3_E_out(clk_3_wires[4]),
    .clk_3_W_in(clk_3_wires[1]),
    .prog_clk_3_E_out(prog_clk_3_wires[4]),
    .prog_clk_3_W_in(prog_clk_3_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[273]),
    .config_enable_E_out(config_enableWires[335]),
    .config_enable_N_out(config_enableWires[334]),
    .config_enable_W_in(config_enableWires[332]),
    .pReset_E_out(pResetWires[335]),
    .pReset_N_out(pResetWires[334]),
    .pReset_W_in(pResetWires[332]),
    .chany_top_in(cby_1__1__65_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__67_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__64_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__58_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__58_ccff_tail),
    .chany_top_out(sb_1__1__45_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__45_ccff_tail)
  );


  sb_1__1_
  sb_7__7_
  (
    .clk_1_N_in(clk_2_wires[98]),
    .clk_1_W_out(clk_1_wires[149]),
    .clk_1_E_out(clk_1_wires[148]),
    .prog_clk_1_N_in(prog_clk_2_wires[98]),
    .prog_clk_1_W_out(prog_clk_1_wires[149]),
    .prog_clk_1_E_out(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[276]),
    .config_enable_E_out(config_enableWires[384]),
    .config_enable_N_out(config_enableWires[383]),
    .config_enable_W_in(config_enableWires[381]),
    .pReset_E_out(pResetWires[384]),
    .pReset_N_out(pResetWires[383]),
    .pReset_W_in(pResetWires[381]),
    .chany_top_in(cby_1__1__66_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__68_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__65_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__59_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__59_ccff_tail),
    .chany_top_out(sb_1__1__46_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__46_ccff_tail)
  );


  sb_1__1_
  sb_7__8_
  (
    .clk_2_S_out(clk_2_wires[97]),
    .clk_2_N_out(clk_2_wires[95]),
    .clk_2_E_in(clk_2_wires[94]),
    .prog_clk_2_S_out(prog_clk_2_wires[97]),
    .prog_clk_2_N_out(prog_clk_2_wires[95]),
    .prog_clk_2_E_in(prog_clk_2_wires[94]),
    .prog_clk_0_N_in(prog_clk_0_wires[279]),
    .config_enable_E_out(config_enableWires[433]),
    .config_enable_N_out(config_enableWires[432]),
    .config_enable_W_in(config_enableWires[430]),
    .pReset_E_out(pResetWires[433]),
    .pReset_N_out(pResetWires[432]),
    .pReset_W_in(pResetWires[430]),
    .chany_top_in(cby_1__1__67_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__69_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__66_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__60_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__60_ccff_tail),
    .chany_top_out(sb_1__1__47_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__47_ccff_tail)
  );


  sb_1__1_
  sb_7__11_
  (
    .clk_1_S_in(clk_2_wires[109]),
    .clk_1_W_out(clk_1_wires[163]),
    .clk_1_E_out(clk_1_wires[162]),
    .prog_clk_1_S_in(prog_clk_2_wires[109]),
    .prog_clk_1_W_out(prog_clk_1_wires[163]),
    .prog_clk_1_E_out(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[288]),
    .config_enable_E_out(config_enableWires[580]),
    .config_enable_N_out(config_enableWires[579]),
    .config_enable_W_in(config_enableWires[577]),
    .pReset_E_out(pResetWires[580]),
    .pReset_N_out(pResetWires[579]),
    .pReset_W_in(pResetWires[577]),
    .chany_top_in(cby_1__1__69_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__71_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__68_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__62_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__62_ccff_tail),
    .chany_top_out(sb_1__1__48_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__48_ccff_tail)
  );


  sb_1__1_
  sb_8__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[296]),
    .config_enable_E_out(config_enableWires[94]),
    .config_enable_N_out(config_enableWires[93]),
    .config_enable_W_in(config_enableWires[91]),
    .pReset_E_out(pResetWires[94]),
    .pReset_N_out(pResetWires[93]),
    .pReset_W_in(pResetWires[91]),
    .chany_top_in(cby_1__1__71_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__72_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__70_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__63_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__63_ccff_tail),
    .chany_top_out(sb_1__1__49_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__49_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__49_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__49_ccff_tail)
  );


  sb_1__1_
  sb_8__4_
  (
    .clk_3_S_out(clk_3_wires[38]),
    .clk_2_N_in(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[33]),
    .clk_2_W_out(clk_2_wires[80]),
    .clk_2_E_out(clk_2_wires[78]),
    .prog_clk_3_S_out(prog_clk_3_wires[38]),
    .prog_clk_2_N_in(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[33]),
    .prog_clk_2_W_out(prog_clk_2_wires[80]),
    .prog_clk_2_E_out(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[305]),
    .config_enable_E_out(config_enableWires[241]),
    .config_enable_N_out(config_enableWires[240]),
    .config_enable_W_in(config_enableWires[238]),
    .pReset_E_out(pResetWires[241]),
    .pReset_N_out(pResetWires[240]),
    .pReset_W_in(pResetWires[238]),
    .chany_top_in(cby_1__1__73_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__74_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__72_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__65_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__65_ccff_tail),
    .chany_top_out(sb_1__1__50_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__50_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__50_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__50_ccff_tail)
  );


  sb_1__1_
  sb_8__5_
  (
    .clk_3_S_out(clk_3_wires[32]),
    .clk_3_N_in(clk_3_wires[29]),
    .prog_clk_3_S_out(prog_clk_3_wires[32]),
    .prog_clk_3_N_in(prog_clk_3_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[308]),
    .config_enable_E_out(config_enableWires[290]),
    .config_enable_N_out(config_enableWires[289]),
    .config_enable_W_in(config_enableWires[287]),
    .pReset_E_out(pResetWires[290]),
    .pReset_N_out(pResetWires[289]),
    .pReset_W_in(pResetWires[287]),
    .chany_top_in(cby_1__1__74_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__75_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__73_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__66_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__66_ccff_tail),
    .chany_top_out(sb_1__1__51_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__51_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__51_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__51_ccff_tail)
  );


  sb_1__1_
  sb_8__6_
  (
    .clk_3_E_out(clk_3_wires[44]),
    .clk_3_S_out(clk_3_wires[28]),
    .clk_3_N_out(clk_3_wires[26]),
    .clk_3_W_in(clk_3_wires[5]),
    .prog_clk_3_E_out(prog_clk_3_wires[44]),
    .prog_clk_3_S_out(prog_clk_3_wires[28]),
    .prog_clk_3_N_out(prog_clk_3_wires[26]),
    .prog_clk_3_W_in(prog_clk_3_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[311]),
    .config_enable_E_out(config_enableWires[339]),
    .config_enable_N_out(config_enableWires[338]),
    .config_enable_W_in(config_enableWires[336]),
    .pReset_E_out(pResetWires[339]),
    .pReset_N_out(pResetWires[338]),
    .pReset_W_in(pResetWires[336]),
    .chany_top_in(cby_1__1__75_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__76_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__74_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__67_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__67_ccff_tail),
    .chany_top_out(sb_1__1__52_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__52_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__52_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__52_ccff_tail)
  );


  sb_1__1_
  sb_8__7_
  (
    .clk_3_N_out(clk_3_wires[30]),
    .clk_3_S_in(clk_3_wires[27]),
    .prog_clk_3_N_out(prog_clk_3_wires[30]),
    .prog_clk_3_S_in(prog_clk_3_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[314]),
    .config_enable_E_out(config_enableWires[388]),
    .config_enable_N_out(config_enableWires[387]),
    .config_enable_W_in(config_enableWires[385]),
    .pReset_E_out(pResetWires[388]),
    .pReset_N_out(pResetWires[387]),
    .pReset_W_in(pResetWires[385]),
    .chany_top_in(cby_1__1__76_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__77_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__75_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__68_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__68_ccff_tail),
    .chany_top_out(sb_1__1__53_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__53_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__53_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__53_ccff_tail)
  );


  sb_1__1_
  sb_8__8_
  (
    .clk_3_N_out(clk_3_wires[36]),
    .clk_2_S_in(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[31]),
    .clk_2_W_out(clk_2_wires[93]),
    .clk_2_E_out(clk_2_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[36]),
    .prog_clk_2_S_in(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[31]),
    .prog_clk_2_W_out(prog_clk_2_wires[93]),
    .prog_clk_2_E_out(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[317]),
    .config_enable_E_out(config_enableWires[437]),
    .config_enable_N_out(config_enableWires[436]),
    .config_enable_W_in(config_enableWires[434]),
    .pReset_E_out(pResetWires[437]),
    .pReset_N_out(pResetWires[436]),
    .pReset_W_in(pResetWires[434]),
    .chany_top_in(cby_1__1__77_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__78_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__76_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__69_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__69_ccff_tail),
    .chany_top_out(sb_1__1__54_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__54_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__54_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__54_ccff_tail)
  );


  sb_1__1_
  sb_8__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[326]),
    .config_enable_E_out(config_enableWires[584]),
    .config_enable_N_out(config_enableWires[583]),
    .config_enable_W_in(config_enableWires[581]),
    .pReset_E_out(pResetWires[584]),
    .pReset_N_out(pResetWires[583]),
    .pReset_W_in(pResetWires[581]),
    .chany_top_in(cby_1__1__79_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__80_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__78_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__71_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__71_ccff_tail),
    .chany_top_out(sb_1__1__55_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__55_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__55_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__55_ccff_tail)
  );


  sb_1__1_
  sb_9__1_
  (
    .clk_1_N_in(clk_2_wires[76]),
    .clk_1_W_out(clk_1_wires[170]),
    .clk_1_E_out(clk_1_wires[169]),
    .prog_clk_1_N_in(prog_clk_2_wires[76]),
    .prog_clk_1_W_out(prog_clk_1_wires[170]),
    .prog_clk_1_E_out(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[334]),
    .config_enable_E_out(config_enableWires[98]),
    .config_enable_N_out(config_enableWires[97]),
    .config_enable_W_in(config_enableWires[95]),
    .pReset_E_out(pResetWires[98]),
    .pReset_N_out(pResetWires[97]),
    .pReset_W_in(pResetWires[95]),
    .chany_top_in(cby_1__1__81_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__81_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__80_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_80_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__72_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_80_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__72_ccff_tail),
    .chany_top_out(sb_1__1__56_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__56_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__56_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__56_ccff_tail)
  );


  sb_1__1_
  sb_9__4_
  (
    .clk_2_S_out(clk_2_wires[88]),
    .clk_2_N_out(clk_2_wires[86]),
    .clk_2_W_in(clk_2_wires[79]),
    .prog_clk_2_S_out(prog_clk_2_wires[88]),
    .prog_clk_2_N_out(prog_clk_2_wires[86]),
    .prog_clk_2_W_in(prog_clk_2_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[343]),
    .config_enable_E_out(config_enableWires[245]),
    .config_enable_N_out(config_enableWires[244]),
    .config_enable_W_in(config_enableWires[242]),
    .pReset_E_out(pResetWires[245]),
    .pReset_N_out(pResetWires[244]),
    .pReset_W_in(pResetWires[242]),
    .chany_top_in(cby_1__1__83_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__83_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__82_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__74_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_82_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__74_ccff_tail),
    .chany_top_out(sb_1__1__57_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__57_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__57_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__57_ccff_tail)
  );


  sb_1__1_
  sb_9__5_
  (
    .clk_1_S_in(clk_2_wires[87]),
    .clk_1_W_out(clk_1_wires[184]),
    .clk_1_E_out(clk_1_wires[183]),
    .prog_clk_1_S_in(prog_clk_2_wires[87]),
    .prog_clk_1_W_out(prog_clk_1_wires[184]),
    .prog_clk_1_E_out(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[346]),
    .config_enable_E_out(config_enableWires[294]),
    .config_enable_N_out(config_enableWires[293]),
    .config_enable_W_in(config_enableWires[291]),
    .pReset_E_out(pResetWires[294]),
    .pReset_N_out(pResetWires[293]),
    .pReset_W_in(pResetWires[291]),
    .chany_top_in(cby_1__1__84_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__84_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__83_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_83_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__75_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_83_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__75_ccff_tail),
    .chany_top_out(sb_1__1__58_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__58_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__58_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__58_ccff_tail)
  );


  sb_1__1_
  sb_9__6_
  (
    .clk_3_E_out(clk_3_wires[48]),
    .clk_3_W_in(clk_3_wires[45]),
    .prog_clk_3_E_out(prog_clk_3_wires[48]),
    .prog_clk_3_W_in(prog_clk_3_wires[45]),
    .prog_clk_0_N_in(prog_clk_0_wires[349]),
    .config_enable_E_out(config_enableWires[343]),
    .config_enable_N_out(config_enableWires[342]),
    .config_enable_W_in(config_enableWires[340]),
    .pReset_E_out(pResetWires[343]),
    .pReset_N_out(pResetWires[342]),
    .pReset_W_in(pResetWires[340]),
    .chany_top_in(cby_1__1__85_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__85_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__84_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_84_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__76_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_84_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__76_ccff_tail),
    .chany_top_out(sb_1__1__59_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__59_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__59_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__59_ccff_tail)
  );


  sb_1__1_
  sb_9__7_
  (
    .clk_1_N_in(clk_2_wires[102]),
    .clk_1_W_out(clk_1_wires[191]),
    .clk_1_E_out(clk_1_wires[190]),
    .prog_clk_1_N_in(prog_clk_2_wires[102]),
    .prog_clk_1_W_out(prog_clk_1_wires[191]),
    .prog_clk_1_E_out(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[352]),
    .config_enable_E_out(config_enableWires[392]),
    .config_enable_N_out(config_enableWires[391]),
    .config_enable_W_in(config_enableWires[389]),
    .pReset_E_out(pResetWires[392]),
    .pReset_N_out(pResetWires[391]),
    .pReset_W_in(pResetWires[389]),
    .chany_top_in(cby_1__1__86_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__86_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__85_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_85_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__77_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_85_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__77_ccff_tail),
    .chany_top_out(sb_1__1__60_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__60_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__60_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__60_ccff_tail)
  );


  sb_1__1_
  sb_9__8_
  (
    .clk_2_S_out(clk_2_wires[101]),
    .clk_2_N_out(clk_2_wires[99]),
    .clk_2_W_in(clk_2_wires[92]),
    .prog_clk_2_S_out(prog_clk_2_wires[101]),
    .prog_clk_2_N_out(prog_clk_2_wires[99]),
    .prog_clk_2_W_in(prog_clk_2_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[355]),
    .config_enable_E_out(config_enableWires[441]),
    .config_enable_N_out(config_enableWires[440]),
    .config_enable_W_in(config_enableWires[438]),
    .pReset_E_out(pResetWires[441]),
    .pReset_N_out(pResetWires[440]),
    .pReset_W_in(pResetWires[438]),
    .chany_top_in(cby_1__1__87_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__87_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__86_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_86_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__78_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_86_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__78_ccff_tail),
    .chany_top_out(sb_1__1__61_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__61_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__61_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__61_ccff_tail)
  );


  sb_1__1_
  sb_9__11_
  (
    .clk_1_S_in(clk_2_wires[111]),
    .clk_1_W_out(clk_1_wires[205]),
    .clk_1_E_out(clk_1_wires[204]),
    .prog_clk_1_S_in(prog_clk_2_wires[111]),
    .prog_clk_1_W_out(prog_clk_1_wires[205]),
    .prog_clk_1_E_out(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[364]),
    .config_enable_E_out(config_enableWires[588]),
    .config_enable_N_out(config_enableWires[587]),
    .config_enable_W_in(config_enableWires[585]),
    .pReset_E_out(pResetWires[588]),
    .pReset_N_out(pResetWires[587]),
    .pReset_W_in(pResetWires[585]),
    .chany_top_in(cby_1__1__89_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__89_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__88_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__80_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_88_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__80_ccff_tail),
    .chany_top_out(sb_1__1__62_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__62_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__62_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__62_ccff_tail)
  );


  sb_1__1_
  sb_10__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[372]),
    .config_enable_E_out(config_enableWires[102]),
    .config_enable_N_out(config_enableWires[101]),
    .config_enable_W_in(config_enableWires[99]),
    .pReset_E_out(pResetWires[102]),
    .pReset_N_out(pResetWires[101]),
    .pReset_W_in(pResetWires[99]),
    .chany_top_in(cby_1__1__91_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__90_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__90_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_90_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__81_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_90_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__81_ccff_tail),
    .chany_top_out(sb_1__1__63_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__63_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__63_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__63_ccff_tail)
  );


  sb_1__1_
  sb_10__4_
  (
    .clk_3_S_out(clk_3_wires[82]),
    .clk_2_N_in(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[77]),
    .clk_2_E_out(clk_2_wires[119]),
    .prog_clk_3_S_out(prog_clk_3_wires[82]),
    .prog_clk_2_N_in(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[77]),
    .prog_clk_2_E_out(prog_clk_2_wires[119]),
    .prog_clk_0_N_in(prog_clk_0_wires[381]),
    .config_enable_E_out(config_enableWires[249]),
    .config_enable_N_out(config_enableWires[248]),
    .config_enable_W_in(config_enableWires[246]),
    .pReset_E_out(pResetWires[249]),
    .pReset_N_out(pResetWires[248]),
    .pReset_W_in(pResetWires[246]),
    .chany_top_in(cby_1__1__93_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__92_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__92_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__83_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_92_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__83_ccff_tail),
    .chany_top_out(sb_1__1__64_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__64_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__64_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__64_ccff_tail)
  );


  sb_1__1_
  sb_10__5_
  (
    .clk_3_S_out(clk_3_wires[76]),
    .clk_3_N_in(clk_3_wires[73]),
    .prog_clk_3_S_out(prog_clk_3_wires[76]),
    .prog_clk_3_N_in(prog_clk_3_wires[73]),
    .prog_clk_0_N_in(prog_clk_0_wires[384]),
    .config_enable_E_out(config_enableWires[298]),
    .config_enable_N_out(config_enableWires[297]),
    .config_enable_W_in(config_enableWires[295]),
    .pReset_E_out(pResetWires[298]),
    .pReset_N_out(pResetWires[297]),
    .pReset_W_in(pResetWires[295]),
    .chany_top_in(cby_1__1__94_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__93_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__93_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_93_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__84_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_93_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__84_ccff_tail),
    .chany_top_out(sb_1__1__65_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__65_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__65_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__65_ccff_tail)
  );


  sb_1__1_
  sb_10__6_
  (
    .clk_3_S_out(clk_3_wires[72]),
    .clk_3_N_out(clk_3_wires[70]),
    .clk_3_W_in(clk_3_wires[49]),
    .prog_clk_3_S_out(prog_clk_3_wires[72]),
    .prog_clk_3_N_out(prog_clk_3_wires[70]),
    .prog_clk_3_W_in(prog_clk_3_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[387]),
    .config_enable_E_out(config_enableWires[347]),
    .config_enable_N_out(config_enableWires[346]),
    .config_enable_W_in(config_enableWires[344]),
    .pReset_E_out(pResetWires[347]),
    .pReset_N_out(pResetWires[346]),
    .pReset_W_in(pResetWires[344]),
    .chany_top_in(cby_1__1__95_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__94_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__94_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_94_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__85_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_94_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__85_ccff_tail),
    .chany_top_out(sb_1__1__66_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__66_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__66_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__66_ccff_tail)
  );


  sb_1__1_
  sb_10__7_
  (
    .clk_3_N_out(clk_3_wires[74]),
    .clk_3_S_in(clk_3_wires[71]),
    .prog_clk_3_N_out(prog_clk_3_wires[74]),
    .prog_clk_3_S_in(prog_clk_3_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[390]),
    .config_enable_E_out(config_enableWires[396]),
    .config_enable_N_out(config_enableWires[395]),
    .config_enable_W_in(config_enableWires[393]),
    .pReset_E_out(pResetWires[396]),
    .pReset_N_out(pResetWires[395]),
    .pReset_W_in(pResetWires[393]),
    .chany_top_in(cby_1__1__96_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__95_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__95_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_95_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__86_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_95_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__86_ccff_tail),
    .chany_top_out(sb_1__1__67_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__67_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__67_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__67_ccff_tail)
  );


  sb_1__1_
  sb_10__8_
  (
    .clk_3_N_out(clk_3_wires[80]),
    .clk_2_S_in(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[75]),
    .clk_2_E_out(clk_2_wires[126]),
    .prog_clk_3_N_out(prog_clk_3_wires[80]),
    .prog_clk_2_S_in(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[75]),
    .prog_clk_2_E_out(prog_clk_2_wires[126]),
    .prog_clk_0_N_in(prog_clk_0_wires[393]),
    .config_enable_E_out(config_enableWires[445]),
    .config_enable_N_out(config_enableWires[444]),
    .config_enable_W_in(config_enableWires[442]),
    .pReset_E_out(pResetWires[445]),
    .pReset_N_out(pResetWires[444]),
    .pReset_W_in(pResetWires[442]),
    .chany_top_in(cby_1__1__97_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__96_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__96_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_96_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__87_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_96_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__87_ccff_tail),
    .chany_top_out(sb_1__1__68_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__68_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__68_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__68_ccff_tail)
  );


  sb_1__1_
  sb_10__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[402]),
    .config_enable_E_out(config_enableWires[592]),
    .config_enable_N_out(config_enableWires[591]),
    .config_enable_W_in(config_enableWires[589]),
    .pReset_E_out(pResetWires[592]),
    .pReset_N_out(pResetWires[591]),
    .pReset_W_in(pResetWires[589]),
    .chany_top_in(cby_1__1__99_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__98_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__98_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__89_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_98_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__89_ccff_tail),
    .chany_top_out(sb_1__1__69_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__69_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__69_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__69_ccff_tail)
  );


  sb_1__1_
  sb_11__1_
  (
    .clk_1_N_in(clk_2_wires[116]),
    .clk_1_W_out(clk_1_wires[212]),
    .clk_1_E_out(clk_1_wires[211]),
    .prog_clk_1_N_in(prog_clk_2_wires[116]),
    .prog_clk_1_W_out(prog_clk_1_wires[212]),
    .prog_clk_1_E_out(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[410]),
    .config_enable_E_out(config_enableWires[106]),
    .config_enable_N_out(config_enableWires[105]),
    .config_enable_W_in(config_enableWires[103]),
    .pReset_E_out(pResetWires[106]),
    .pReset_N_out(pResetWires[105]),
    .pReset_W_in(pResetWires[103]),
    .chany_top_in(cby_1__1__101_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__99_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__100_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_100_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__90_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_100_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__90_ccff_tail),
    .chany_top_out(sb_1__1__70_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__70_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__70_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__70_ccff_tail)
  );


  sb_1__1_
  sb_11__4_
  (
    .clk_2_S_out(clk_2_wires[122]),
    .clk_2_N_out(clk_2_wires[120]),
    .clk_2_W_in(clk_2_wires[118]),
    .prog_clk_2_S_out(prog_clk_2_wires[122]),
    .prog_clk_2_N_out(prog_clk_2_wires[120]),
    .prog_clk_2_W_in(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[419]),
    .config_enable_E_out(config_enableWires[253]),
    .config_enable_N_out(config_enableWires[252]),
    .config_enable_W_in(config_enableWires[250]),
    .pReset_E_out(pResetWires[253]),
    .pReset_N_out(pResetWires[252]),
    .pReset_W_in(pResetWires[250]),
    .chany_top_in(cby_1__1__103_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__101_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__102_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__92_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_102_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__92_ccff_tail),
    .chany_top_out(sb_1__1__71_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__71_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__71_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__71_ccff_tail)
  );


  sb_1__1_
  sb_11__5_
  (
    .clk_1_S_in(clk_2_wires[121]),
    .clk_1_W_out(clk_1_wires[226]),
    .clk_1_E_out(clk_1_wires[225]),
    .prog_clk_1_S_in(prog_clk_2_wires[121]),
    .prog_clk_1_W_out(prog_clk_1_wires[226]),
    .prog_clk_1_E_out(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[422]),
    .config_enable_E_out(config_enableWires[302]),
    .config_enable_N_out(config_enableWires[301]),
    .config_enable_W_in(config_enableWires[299]),
    .pReset_E_out(pResetWires[302]),
    .pReset_N_out(pResetWires[301]),
    .pReset_W_in(pResetWires[299]),
    .chany_top_in(cby_1__1__104_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__102_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__103_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_103_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__93_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_103_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__93_ccff_tail),
    .chany_top_out(sb_1__1__72_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__72_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__72_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__72_ccff_tail)
  );


  sb_1__1_
  sb_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[425]),
    .config_enable_E_out(config_enableWires[351]),
    .config_enable_N_out(config_enableWires[350]),
    .config_enable_W_in(config_enableWires[348]),
    .pReset_E_out(pResetWires[351]),
    .pReset_N_out(pResetWires[350]),
    .pReset_W_in(pResetWires[348]),
    .chany_top_in(cby_1__1__105_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__103_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__104_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_104_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__94_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_104_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__94_ccff_tail),
    .chany_top_out(sb_1__1__73_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__73_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__73_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__73_ccff_tail)
  );


  sb_1__1_
  sb_11__7_
  (
    .clk_1_N_in(clk_2_wires[130]),
    .clk_1_W_out(clk_1_wires[233]),
    .clk_1_E_out(clk_1_wires[232]),
    .prog_clk_1_N_in(prog_clk_2_wires[130]),
    .prog_clk_1_W_out(prog_clk_1_wires[233]),
    .prog_clk_1_E_out(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[428]),
    .config_enable_E_out(config_enableWires[400]),
    .config_enable_N_out(config_enableWires[399]),
    .config_enable_W_in(config_enableWires[397]),
    .pReset_E_out(pResetWires[400]),
    .pReset_N_out(pResetWires[399]),
    .pReset_W_in(pResetWires[397]),
    .chany_top_in(cby_1__1__106_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__104_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__105_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_105_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__95_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_105_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__95_ccff_tail),
    .chany_top_out(sb_1__1__74_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__74_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__74_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__74_ccff_tail)
  );


  sb_1__1_
  sb_11__8_
  (
    .clk_2_S_out(clk_2_wires[129]),
    .clk_2_N_out(clk_2_wires[127]),
    .clk_2_W_in(clk_2_wires[125]),
    .prog_clk_2_S_out(prog_clk_2_wires[129]),
    .prog_clk_2_N_out(prog_clk_2_wires[127]),
    .prog_clk_2_W_in(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[431]),
    .config_enable_E_out(config_enableWires[449]),
    .config_enable_N_out(config_enableWires[448]),
    .config_enable_W_in(config_enableWires[446]),
    .pReset_E_out(pResetWires[449]),
    .pReset_N_out(pResetWires[448]),
    .pReset_W_in(pResetWires[446]),
    .chany_top_in(cby_1__1__107_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__105_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__106_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_106_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__96_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_106_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__96_ccff_tail),
    .chany_top_out(sb_1__1__75_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__75_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__75_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__75_ccff_tail)
  );


  sb_1__1_
  sb_11__11_
  (
    .clk_1_S_in(clk_2_wires[135]),
    .clk_1_W_out(clk_1_wires[247]),
    .clk_1_E_out(clk_1_wires[246]),
    .prog_clk_1_S_in(prog_clk_2_wires[135]),
    .prog_clk_1_W_out(prog_clk_1_wires[247]),
    .prog_clk_1_E_out(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[440]),
    .config_enable_E_out(config_enableWires[596]),
    .config_enable_N_out(config_enableWires[595]),
    .config_enable_W_in(config_enableWires[593]),
    .pReset_E_out(pResetWires[596]),
    .pReset_N_out(pResetWires[595]),
    .pReset_W_in(pResetWires[593]),
    .chany_top_in(cby_1__1__109_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__1__107_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__108_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__98_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_108_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__98_ccff_tail),
    .chany_top_out(sb_1__1__76_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__76_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__76_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__76_ccff_tail)
  );


  sb_1__2_
  sb_1__2_
  (
    .clk_2_S_out(clk_2_wires[3]),
    .clk_2_E_in(clk_2_wires[1]),
    .prog_clk_2_S_out(prog_clk_2_wires[3]),
    .prog_clk_2_E_in(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[13]),
    .config_enable_E_in(config_enableWires[115]),
    .config_enable_N_out(config_enableWires[114]),
    .config_enable_W_out(config_enableWires[111]),
    .pReset_E_in(pResetWires[115]),
    .pReset_N_out(pResetWires[114]),
    .pReset_W_out(pResetWires[111]),
    .chany_top_in(cby_1__3__0_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__1_ccff_tail),
    .chany_top_out(sb_1__2__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__0_ccff_tail)
  );


  sb_1__2_
  sb_1__9_
  (
    .clk_1_S_in(clk_2_wires[16]),
    .clk_1_W_out(clk_1_wires[30]),
    .clk_1_E_out(clk_1_wires[29]),
    .prog_clk_1_S_in(prog_clk_2_wires[16]),
    .prog_clk_1_W_out(prog_clk_1_wires[30]),
    .prog_clk_1_E_out(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[48]),
    .config_enable_E_in(config_enableWires[458]),
    .config_enable_N_out(config_enableWires[457]),
    .config_enable_W_out(config_enableWires[454]),
    .pReset_E_in(pResetWires[458]),
    .pReset_N_out(pResetWires[457]),
    .pReset_W_out(pResetWires[454]),
    .chany_top_in(cby_1__3__1_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__7_ccff_tail),
    .chany_top_out(sb_1__2__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__1_ccff_tail)
  );


  sb_1__2_
  sb_3__2_
  (
    .clk_2_S_out(clk_2_wires[29]),
    .clk_2_E_in(clk_2_wires[28]),
    .prog_clk_2_S_out(prog_clk_2_wires[29]),
    .prog_clk_2_E_in(prog_clk_2_wires[28]),
    .prog_clk_0_N_in(prog_clk_0_wires[109]),
    .config_enable_E_in(config_enableWires[123]),
    .config_enable_N_out(config_enableWires[122]),
    .config_enable_W_out(config_enableWires[120]),
    .pReset_E_in(pResetWires[123]),
    .pReset_N_out(pResetWires[122]),
    .pReset_W_out(pResetWires[120]),
    .chany_top_in(cby_1__3__2_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__19_ccff_tail),
    .chany_top_out(sb_1__2__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__2_ccff_tail)
  );


  sb_1__2_
  sb_3__9_
  (
    .clk_1_S_in(clk_2_wires[52]),
    .clk_1_W_out(clk_1_wires[72]),
    .clk_1_E_out(clk_1_wires[71]),
    .prog_clk_1_S_in(prog_clk_2_wires[52]),
    .prog_clk_1_W_out(prog_clk_1_wires[72]),
    .prog_clk_1_E_out(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[130]),
    .config_enable_E_in(config_enableWires[466]),
    .config_enable_N_out(config_enableWires[465]),
    .config_enable_W_out(config_enableWires[463]),
    .pReset_E_in(pResetWires[466]),
    .pReset_N_out(pResetWires[465]),
    .pReset_W_out(pResetWires[463]),
    .chany_top_in(cby_1__3__3_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__25_ccff_tail),
    .chany_top_out(sb_1__2__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__3_ccff_tail)
  );


  sb_1__2_
  sb_5__2_
  (
    .clk_2_S_out(clk_2_wires[31]),
    .clk_2_W_in(clk_2_wires[26]),
    .prog_clk_2_S_out(prog_clk_2_wires[31]),
    .prog_clk_2_W_in(prog_clk_2_wires[26]),
    .prog_clk_0_N_in(prog_clk_0_wires[185]),
    .config_enable_E_in(config_enableWires[131]),
    .config_enable_N_out(config_enableWires[130]),
    .config_enable_W_out(config_enableWires[128]),
    .pReset_E_in(pResetWires[131]),
    .pReset_N_out(pResetWires[130]),
    .pReset_W_out(pResetWires[128]),
    .chany_top_in(cby_1__3__4_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__37_ccff_tail),
    .chany_top_out(sb_1__2__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__4_ccff_tail)
  );


  sb_1__2_
  sb_5__9_
  (
    .clk_1_S_in(clk_2_wires[56]),
    .clk_1_W_out(clk_1_wires[114]),
    .clk_1_E_out(clk_1_wires[113]),
    .prog_clk_1_S_in(prog_clk_2_wires[56]),
    .prog_clk_1_W_out(prog_clk_1_wires[114]),
    .prog_clk_1_E_out(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[206]),
    .config_enable_E_in(config_enableWires[474]),
    .config_enable_N_out(config_enableWires[473]),
    .config_enable_W_out(config_enableWires[471]),
    .pReset_E_in(pResetWires[474]),
    .pReset_N_out(pResetWires[473]),
    .pReset_W_out(pResetWires[471]),
    .chany_top_in(cby_1__3__5_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__43_ccff_tail),
    .chany_top_out(sb_1__2__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__5_ccff_tail)
  );


  sb_1__2_
  sb_7__2_
  (
    .clk_2_S_out(clk_2_wires[73]),
    .clk_2_E_in(clk_2_wires[72]),
    .prog_clk_2_S_out(prog_clk_2_wires[73]),
    .prog_clk_2_E_in(prog_clk_2_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[261]),
    .config_enable_E_out(config_enableWires[139]),
    .config_enable_N_out(config_enableWires[138]),
    .config_enable_W_in(config_enableWires[136]),
    .pReset_E_out(pResetWires[139]),
    .pReset_N_out(pResetWires[138]),
    .pReset_W_in(pResetWires[136]),
    .chany_top_in(cby_1__3__6_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__64_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__61_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__55_ccff_tail),
    .chany_top_out(sb_1__2__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__6_ccff_tail)
  );


  sb_1__2_
  sb_7__9_
  (
    .clk_1_S_in(clk_2_wires[96]),
    .clk_1_W_out(clk_1_wires[156]),
    .clk_1_E_out(clk_1_wires[155]),
    .prog_clk_1_S_in(prog_clk_2_wires[96]),
    .prog_clk_1_W_out(prog_clk_1_wires[156]),
    .prog_clk_1_E_out(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[282]),
    .config_enable_E_out(config_enableWires[482]),
    .config_enable_N_out(config_enableWires[481]),
    .config_enable_W_in(config_enableWires[479]),
    .pReset_E_out(pResetWires[482]),
    .pReset_N_out(pResetWires[481]),
    .pReset_W_in(pResetWires[479]),
    .chany_top_in(cby_1__3__7_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__70_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__67_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__61_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__61_ccff_tail),
    .chany_top_out(sb_1__2__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__7_ccff_tail)
  );


  sb_1__2_
  sb_9__2_
  (
    .clk_2_S_out(clk_2_wires[75]),
    .clk_2_W_in(clk_2_wires[70]),
    .prog_clk_2_S_out(prog_clk_2_wires[75]),
    .prog_clk_2_W_in(prog_clk_2_wires[70]),
    .prog_clk_0_N_in(prog_clk_0_wires[337]),
    .config_enable_E_out(config_enableWires[147]),
    .config_enable_N_out(config_enableWires[146]),
    .config_enable_W_in(config_enableWires[144]),
    .pReset_E_out(pResetWires[147]),
    .pReset_N_out(pResetWires[146]),
    .pReset_W_in(pResetWires[144]),
    .chany_top_in(cby_1__3__8_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__82_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__81_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_81_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__73_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__73_ccff_tail),
    .chany_top_out(sb_1__2__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__8_ccff_tail)
  );


  sb_1__2_
  sb_9__9_
  (
    .clk_1_S_in(clk_2_wires[100]),
    .clk_1_W_out(clk_1_wires[198]),
    .clk_1_E_out(clk_1_wires[197]),
    .prog_clk_1_S_in(prog_clk_2_wires[100]),
    .prog_clk_1_W_out(prog_clk_1_wires[198]),
    .prog_clk_1_E_out(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[358]),
    .config_enable_E_out(config_enableWires[490]),
    .config_enable_N_out(config_enableWires[489]),
    .config_enable_W_in(config_enableWires[487]),
    .pReset_E_out(pResetWires[490]),
    .pReset_N_out(pResetWires[489]),
    .pReset_W_in(pResetWires[487]),
    .chany_top_in(cby_1__3__9_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__88_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__87_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_87_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__79_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__79_ccff_tail),
    .chany_top_out(sb_1__2__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__9_ccff_tail)
  );


  sb_1__2_
  sb_11__2_
  (
    .clk_2_S_out(clk_2_wires[115]),
    .clk_2_W_in(clk_2_wires[113]),
    .prog_clk_2_S_out(prog_clk_2_wires[115]),
    .prog_clk_2_W_in(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[413]),
    .config_enable_E_out(config_enableWires[155]),
    .config_enable_N_out(config_enableWires[154]),
    .config_enable_W_in(config_enableWires[152]),
    .pReset_E_out(pResetWires[155]),
    .pReset_N_out(pResetWires[154]),
    .pReset_W_in(pResetWires[152]),
    .chany_top_in(cby_1__3__10_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__100_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__101_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_101_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__91_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__91_ccff_tail),
    .chany_top_out(sb_1__2__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__10_ccff_tail)
  );


  sb_1__2_
  sb_11__9_
  (
    .clk_1_S_in(clk_2_wires[128]),
    .clk_1_W_out(clk_1_wires[240]),
    .clk_1_E_out(clk_1_wires[239]),
    .prog_clk_1_S_in(prog_clk_2_wires[128]),
    .prog_clk_1_W_out(prog_clk_1_wires[240]),
    .prog_clk_1_E_out(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[434]),
    .config_enable_E_out(config_enableWires[498]),
    .config_enable_N_out(config_enableWires[497]),
    .config_enable_W_in(config_enableWires[495]),
    .pReset_E_out(pResetWires[498]),
    .pReset_N_out(pResetWires[497]),
    .pReset_W_in(pResetWires[495]),
    .chany_top_in(cby_1__3__11_chany_bottom_out[0:19]),
    .chanx_right_in(cbx_1__1__106_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__107_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_107_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__97_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__97_ccff_tail),
    .chany_top_out(sb_1__2__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__2__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__2__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__2__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__2__11_ccff_tail)
  );


  sb_1__3_
  sb_1__3_
  (
    .clk_1_N_in(clk_2_wires[11]),
    .clk_1_W_out(clk_1_wires[9]),
    .clk_1_E_out(clk_1_wires[8]),
    .prog_clk_1_N_in(prog_clk_2_wires[11]),
    .prog_clk_1_W_out(prog_clk_1_wires[9]),
    .prog_clk_1_E_out(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[18]),
    .config_enable_E_in(config_enableWires[164]),
    .config_enable_N_out(config_enableWires[163]),
    .config_enable_W_out(config_enableWires[160]),
    .pReset_E_in(pResetWires[164]),
    .pReset_N_out(pResetWires[163]),
    .pReset_W_out(pResetWires[160]),
    .chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__0_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__0_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_0_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__0_ccff_tail),
    .chany_top_out(sb_1__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__0_ccff_tail)
  );


  sb_1__3_
  sb_1__10_
  (
    .clk_2_N_out(clk_2_wires[22]),
    .clk_2_E_in(clk_2_wires[20]),
    .prog_clk_2_N_out(prog_clk_2_wires[22]),
    .prog_clk_2_E_in(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[53]),
    .config_enable_E_in(config_enableWires[507]),
    .config_enable_N_out(config_enableWires[506]),
    .config_enable_W_out(config_enableWires[503]),
    .pReset_E_in(pResetWires[507]),
    .pReset_N_out(pResetWires[506]),
    .pReset_W_out(pResetWires[503]),
    .chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__1_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__1_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_1_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__1_ccff_tail),
    .chany_top_out(sb_1__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__1_ccff_tail)
  );


  sb_1__3_
  sb_3__3_
  (
    .clk_1_N_in(clk_2_wires[41]),
    .clk_1_W_out(clk_1_wires[51]),
    .clk_1_E_out(clk_1_wires[50]),
    .prog_clk_1_N_in(prog_clk_2_wires[41]),
    .prog_clk_1_W_out(prog_clk_1_wires[51]),
    .prog_clk_1_E_out(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[112]),
    .config_enable_E_in(config_enableWires[172]),
    .config_enable_N_out(config_enableWires[171]),
    .config_enable_W_out(config_enableWires[169]),
    .pReset_E_in(pResetWires[172]),
    .pReset_N_out(pResetWires[171]),
    .pReset_W_out(pResetWires[169]),
    .chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__2_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__2_ccff_tail),
    .chany_top_out(sb_1__3__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__2_ccff_tail)
  );


  sb_1__3_
  sb_3__10_
  (
    .clk_2_N_out(clk_2_wires[64]),
    .clk_2_E_in(clk_2_wires[63]),
    .prog_clk_2_N_out(prog_clk_2_wires[64]),
    .prog_clk_2_E_in(prog_clk_2_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[133]),
    .config_enable_E_in(config_enableWires[515]),
    .config_enable_N_out(config_enableWires[514]),
    .config_enable_W_out(config_enableWires[512]),
    .pReset_E_in(pResetWires[515]),
    .pReset_N_out(pResetWires[514]),
    .pReset_W_out(pResetWires[512]),
    .chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__3_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__3_ccff_tail),
    .chany_top_out(sb_1__3__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__3_ccff_tail)
  );


  sb_1__3_
  sb_5__3_
  (
    .clk_1_N_in(clk_2_wires[45]),
    .clk_1_W_out(clk_1_wires[93]),
    .clk_1_E_out(clk_1_wires[92]),
    .prog_clk_1_N_in(prog_clk_2_wires[45]),
    .prog_clk_1_W_out(prog_clk_1_wires[93]),
    .prog_clk_1_E_out(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[188]),
    .config_enable_E_in(config_enableWires[180]),
    .config_enable_N_out(config_enableWires[179]),
    .config_enable_W_out(config_enableWires[177]),
    .pReset_E_in(pResetWires[180]),
    .pReset_N_out(pResetWires[179]),
    .pReset_W_out(pResetWires[177]),
    .chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__4_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__4_ccff_tail),
    .chany_top_out(sb_1__3__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__4_ccff_tail)
  );


  sb_1__3_
  sb_5__10_
  (
    .clk_2_N_out(clk_2_wires[66]),
    .clk_2_W_in(clk_2_wires[61]),
    .prog_clk_2_N_out(prog_clk_2_wires[66]),
    .prog_clk_2_W_in(prog_clk_2_wires[61]),
    .prog_clk_0_N_in(prog_clk_0_wires[209]),
    .config_enable_E_in(config_enableWires[523]),
    .config_enable_N_out(config_enableWires[522]),
    .config_enable_W_out(config_enableWires[520]),
    .pReset_E_in(pResetWires[523]),
    .pReset_N_out(pResetWires[522]),
    .pReset_W_out(pResetWires[520]),
    .chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__5_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__5_ccff_tail),
    .chany_top_out(sb_1__3__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__5_ccff_tail)
  );


  sb_1__3_
  sb_7__3_
  (
    .clk_1_N_in(clk_2_wires[85]),
    .clk_1_W_out(clk_1_wires[135]),
    .clk_1_E_out(clk_1_wires[134]),
    .prog_clk_1_N_in(prog_clk_2_wires[85]),
    .prog_clk_1_W_out(prog_clk_1_wires[135]),
    .prog_clk_1_E_out(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[264]),
    .config_enable_E_out(config_enableWires[188]),
    .config_enable_N_out(config_enableWires[187]),
    .config_enable_W_in(config_enableWires[185]),
    .pReset_E_out(pResetWires[188]),
    .pReset_N_out(pResetWires[187]),
    .pReset_W_in(pResetWires[185]),
    .chany_top_in(cby_1__1__62_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__6_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__6_ccff_tail),
    .chany_top_out(sb_1__3__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__6_ccff_tail)
  );


  sb_1__3_
  sb_7__10_
  (
    .clk_2_N_out(clk_2_wires[108]),
    .clk_2_E_in(clk_2_wires[107]),
    .prog_clk_2_N_out(prog_clk_2_wires[108]),
    .prog_clk_2_E_in(prog_clk_2_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[285]),
    .config_enable_E_out(config_enableWires[531]),
    .config_enable_N_out(config_enableWires[530]),
    .config_enable_W_in(config_enableWires[528]),
    .pReset_E_out(pResetWires[531]),
    .pReset_N_out(pResetWires[530]),
    .pReset_W_in(pResetWires[528]),
    .chany_top_in(cby_1__1__68_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__7_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__7_ccff_tail),
    .chany_top_out(sb_1__3__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__7_ccff_tail)
  );


  sb_1__3_
  sb_9__3_
  (
    .clk_1_N_in(clk_2_wires[89]),
    .clk_1_W_out(clk_1_wires[177]),
    .clk_1_E_out(clk_1_wires[176]),
    .prog_clk_1_N_in(prog_clk_2_wires[89]),
    .prog_clk_1_W_out(prog_clk_1_wires[177]),
    .prog_clk_1_E_out(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[340]),
    .config_enable_E_out(config_enableWires[196]),
    .config_enable_N_out(config_enableWires[195]),
    .config_enable_W_in(config_enableWires[193]),
    .pReset_E_out(pResetWires[196]),
    .pReset_N_out(pResetWires[195]),
    .pReset_W_in(pResetWires[193]),
    .chany_top_in(cby_1__1__82_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_82_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__8_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__8_ccff_tail),
    .chany_top_out(sb_1__3__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__8_ccff_tail)
  );


  sb_1__3_
  sb_9__10_
  (
    .clk_2_N_out(clk_2_wires[110]),
    .clk_2_W_in(clk_2_wires[105]),
    .prog_clk_2_N_out(prog_clk_2_wires[110]),
    .prog_clk_2_W_in(prog_clk_2_wires[105]),
    .prog_clk_0_N_in(prog_clk_0_wires[361]),
    .config_enable_E_out(config_enableWires[539]),
    .config_enable_N_out(config_enableWires[538]),
    .config_enable_W_in(config_enableWires[536]),
    .pReset_E_out(pResetWires[539]),
    .pReset_N_out(pResetWires[538]),
    .pReset_W_in(pResetWires[536]),
    .chany_top_in(cby_1__1__88_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_88_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__9_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__9_ccff_tail),
    .chany_top_out(sb_1__3__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__9_ccff_tail)
  );


  sb_1__3_
  sb_11__3_
  (
    .clk_1_N_in(clk_2_wires[123]),
    .clk_1_W_out(clk_1_wires[219]),
    .clk_1_E_out(clk_1_wires[218]),
    .prog_clk_1_N_in(prog_clk_2_wires[123]),
    .prog_clk_1_W_out(prog_clk_1_wires[219]),
    .prog_clk_1_E_out(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[416]),
    .config_enable_E_out(config_enableWires[204]),
    .config_enable_N_out(config_enableWires[203]),
    .config_enable_W_in(config_enableWires[201]),
    .pReset_E_out(pResetWires[204]),
    .pReset_N_out(pResetWires[203]),
    .pReset_W_in(pResetWires[201]),
    .chany_top_in(cby_1__1__102_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_102_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__10_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__10_ccff_tail),
    .chany_top_out(sb_1__3__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__10_ccff_tail)
  );


  sb_1__3_
  sb_11__10_
  (
    .clk_2_N_out(clk_2_wires[134]),
    .clk_2_W_in(clk_2_wires[132]),
    .prog_clk_2_N_out(prog_clk_2_wires[134]),
    .prog_clk_2_W_in(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[437]),
    .config_enable_E_out(config_enableWires[547]),
    .config_enable_N_out(config_enableWires[546]),
    .config_enable_W_in(config_enableWires[544]),
    .pReset_E_out(pResetWires[547]),
    .pReset_N_out(pResetWires[546]),
    .pReset_W_in(pResetWires[544]),
    .chany_top_in(cby_1__1__108_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_108_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_2__3__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_upper),
    .right_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_upper),
    .chany_bottom_in(cby_1__3__11_chany_top_out[0:19]),
    .chanx_left_in(cbx_1__3__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_lower),
    .ccff_head(cbx_1__3__11_ccff_tail),
    .chany_top_out(sb_1__3__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__3__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__3__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__3__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__3__11_ccff_tail)
  );


  sb_1__4_
  sb_1__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[60]),
    .config_enable_E_in(config_enableWires[604]),
    .config_enable_W_out(config_enableWires[601]),
    .pReset_E_in(pResetWires[604]),
    .pReset_W_out(pResetWires[601]),
    .chanx_right_in(cbx_1__12__1_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__0_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_1_ccff_tail),
    .chanx_right_out(sb_1__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__0_ccff_tail)
  );


  sb_1__4_
  sb_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[100]),
    .config_enable_E_in(config_enableWires[607]),
    .config_enable_W_out(config_enableWires[605]),
    .sc_head_E_out(sc_headWires[53]),
    .sc_head_W_in(sc_headWires[52]),
    .pReset_E_in(pResetWires[607]),
    .pReset_W_out(pResetWires[605]),
    .chanx_right_in(cbx_1__12__2_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__1_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_2_ccff_tail),
    .chanx_right_out(sb_1__12__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__1_ccff_tail)
  );


  sb_1__4_
  sb_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[138]),
    .config_enable_E_in(config_enableWires[610]),
    .config_enable_W_out(config_enableWires[608]),
    .pReset_E_in(pResetWires[610]),
    .pReset_W_out(pResetWires[608]),
    .chanx_right_in(cbx_1__12__3_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__2_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_3_ccff_tail),
    .chanx_right_out(sb_1__12__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__2_ccff_tail)
  );


  sb_1__4_
  sb_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[176]),
    .config_enable_E_in(config_enableWires[613]),
    .config_enable_W_out(config_enableWires[611]),
    .sc_head_E_out(sc_headWires[105]),
    .sc_head_W_in(sc_headWires[104]),
    .pReset_E_in(pResetWires[613]),
    .pReset_W_out(pResetWires[611]),
    .chanx_right_in(cbx_1__12__4_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__3_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_4_ccff_tail),
    .chanx_right_out(sb_1__12__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__3_ccff_tail)
  );


  sb_1__4_
  sb_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[214]),
    .config_enable_E_in(config_enableWires[616]),
    .config_enable_W_out(config_enableWires[614]),
    .pReset_E_in(pResetWires[616]),
    .pReset_W_out(pResetWires[614]),
    .chanx_right_in(cbx_1__12__5_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__4_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_5_ccff_tail),
    .chanx_right_out(sb_1__12__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__4_ccff_tail)
  );


  sb_1__4_
  sb_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[252]),
    .config_enable_E_out(config_enableWires[619]),
    .config_enable_W_out(config_enableWires[617]),
    .config_enable_S_in(config_enableWires[24]),
    .sc_head_E_out(sc_headWires[157]),
    .sc_head_W_in(sc_headWires[156]),
    .pReset_E_out(pResetWires[619]),
    .pReset_W_out(pResetWires[617]),
    .pReset_S_in(pResetWires[24]),
    .chanx_right_in(cbx_1__12__6_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__59_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__5_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_6_ccff_tail),
    .chanx_right_out(sb_1__12__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__5_ccff_tail)
  );


  sb_1__4_
  sb_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[290]),
    .config_enable_E_out(config_enableWires[622]),
    .config_enable_W_in(config_enableWires[620]),
    .pReset_E_out(pResetWires[622]),
    .pReset_W_in(pResetWires[620]),
    .chanx_right_in(cbx_1__12__7_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__69_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__6_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_7_ccff_tail),
    .chanx_right_out(sb_1__12__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__6_ccff_tail)
  );


  sb_1__4_
  sb_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[328]),
    .config_enable_E_out(config_enableWires[625]),
    .config_enable_W_in(config_enableWires[623]),
    .sc_head_E_out(sc_headWires[209]),
    .sc_head_W_in(sc_headWires[208]),
    .pReset_E_out(pResetWires[625]),
    .pReset_W_in(pResetWires[623]),
    .chanx_right_in(cbx_1__12__8_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__79_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__7_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_8_ccff_tail),
    .chanx_right_out(sb_1__12__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__7_ccff_tail)
  );


  sb_1__4_
  sb_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[366]),
    .config_enable_E_out(config_enableWires[628]),
    .config_enable_W_in(config_enableWires[626]),
    .pReset_E_out(pResetWires[628]),
    .pReset_W_in(pResetWires[626]),
    .chanx_right_in(cbx_1__12__9_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__89_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_89_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__8_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_89_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_9_ccff_tail),
    .chanx_right_out(sb_1__12__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__8_ccff_tail)
  );


  sb_1__4_
  sb_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[404]),
    .config_enable_E_out(config_enableWires[631]),
    .config_enable_W_in(config_enableWires[629]),
    .sc_head_E_out(sc_headWires[261]),
    .sc_head_W_in(sc_headWires[260]),
    .pReset_E_out(pResetWires[631]),
    .pReset_W_in(pResetWires[629]),
    .chanx_right_in(cbx_1__12__10_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__99_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_99_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__9_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_99_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_10_ccff_tail),
    .chanx_right_out(sb_1__12__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__9_ccff_tail)
  );


  sb_1__4_
  sb_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[442]),
    .config_enable_E_out(config_enableWires[634]),
    .config_enable_W_in(config_enableWires[632]),
    .pReset_E_out(pResetWires[634]),
    .pReset_W_in(pResetWires[632]),
    .chanx_right_in(cbx_1__12__11_chanx_left_out[0:19]),
    .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__109_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_109_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__10_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_109_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(grid_io_top_top_11_ccff_tail),
    .chanx_right_out(sb_1__12__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__10_ccff_tail)
  );


  sb_2__2_
  sb_2__2_
  (
    .clk_2_N_in(clk_3_wires[69]),
    .clk_2_W_out(clk_2_wires[2]),
    .prog_clk_2_N_in(prog_clk_3_wires[69]),
    .prog_clk_2_W_out(prog_clk_2_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[71]),
    .config_enable_E_in(config_enableWires[119]),
    .config_enable_N_out(config_enableWires[118]),
    .config_enable_W_out(config_enableWires[116]),
    .pReset_E_in(pResetWires[119]),
    .pReset_N_out(pResetWires[118]),
    .pReset_W_out(pResetWires[116]),
    .chany_top_in(cby_2__3__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__10_ccff_tail),
    .chany_top_out(sb_2__2__0_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__0_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__0_ccff_tail)
  );


  sb_2__2_
  sb_2__9_
  (
    .clk_3_N_out(clk_3_wires[66]),
    .clk_3_S_in(clk_3_wires[63]),
    .prog_clk_3_N_out(prog_clk_3_wires[66]),
    .prog_clk_3_S_in(prog_clk_3_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[92]),
    .config_enable_E_in(config_enableWires[462]),
    .config_enable_N_out(config_enableWires[461]),
    .config_enable_W_out(config_enableWires[459]),
    .pReset_E_in(pResetWires[462]),
    .pReset_N_out(pResetWires[461]),
    .pReset_W_out(pResetWires[459]),
    .chany_top_in(cby_2__3__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__16_ccff_tail),
    .chany_top_out(sb_2__2__1_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__1_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__1_ccff_tail)
  );


  sb_2__2_
  sb_4__2_
  (
    .clk_2_N_in(clk_3_wires[25]),
    .clk_2_W_out(clk_2_wires[27]),
    .clk_2_E_out(clk_2_wires[25]),
    .prog_clk_2_N_in(prog_clk_3_wires[25]),
    .prog_clk_2_W_out(prog_clk_2_wires[27]),
    .prog_clk_2_E_out(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[147]),
    .config_enable_E_in(config_enableWires[127]),
    .config_enable_N_out(config_enableWires[126]),
    .config_enable_W_out(config_enableWires[124]),
    .pReset_E_in(pResetWires[127]),
    .pReset_N_out(pResetWires[126]),
    .pReset_W_out(pResetWires[124]),
    .chany_top_in(cby_2__3__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__28_ccff_tail),
    .chany_top_out(sb_2__2__2_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__2_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__2_ccff_tail)
  );


  sb_2__2_
  sb_4__9_
  (
    .clk_3_N_out(clk_3_wires[22]),
    .clk_3_S_in(clk_3_wires[19]),
    .prog_clk_3_N_out(prog_clk_3_wires[22]),
    .prog_clk_3_S_in(prog_clk_3_wires[19]),
    .prog_clk_0_N_in(prog_clk_0_wires[168]),
    .config_enable_E_in(config_enableWires[470]),
    .config_enable_N_out(config_enableWires[469]),
    .config_enable_W_out(config_enableWires[467]),
    .pReset_E_in(pResetWires[470]),
    .pReset_N_out(pResetWires[469]),
    .pReset_W_out(pResetWires[467]),
    .chany_top_in(cby_2__3__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__34_ccff_tail),
    .chany_top_out(sb_2__2__3_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__3_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__3_ccff_tail)
  );


  sb_2__2_
  sb_6__2_
  (
    .clk_3_N_out(clk_3_wires[94]),
    .clk_3_S_in(clk_3_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[94]),
    .prog_clk_3_S_in(prog_clk_3_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[223]),
    .config_enable_E_out(config_enableWires[135]),
    .config_enable_W_out(config_enableWires[132]),
    .config_enable_N_out(config_enableWires[134]),
    .config_enable_S_in(config_enableWires[4]),
    .reset_N_out(resetWires[5]),
    .reset_S_in(resetWires[4]),
    .Test_en_N_out(Test_enWires[5]),
    .Test_en_S_in(Test_enWires[4]),
    .pReset_E_out(pResetWires[135]),
    .pReset_W_out(pResetWires[132]),
    .pReset_N_out(pResetWires[134]),
    .pReset_S_in(pResetWires[4]),
    .chany_top_in(cby_2__3__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__46_ccff_tail),
    .chany_top_out(sb_2__2__4_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__4_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__4_ccff_tail)
  );


  sb_2__2_
  sb_6__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[244]),
    .config_enable_E_out(config_enableWires[478]),
    .config_enable_W_out(config_enableWires[475]),
    .config_enable_N_out(config_enableWires[477]),
    .config_enable_S_in(config_enableWires[18]),
    .reset_N_out(resetWires[19]),
    .reset_S_in(resetWires[18]),
    .Test_en_N_out(Test_enWires[19]),
    .Test_en_S_in(Test_enWires[18]),
    .pReset_E_out(pResetWires[478]),
    .pReset_W_out(pResetWires[475]),
    .pReset_N_out(pResetWires[477]),
    .pReset_S_in(pResetWires[18]),
    .chany_top_in(cby_2__3__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__61_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__57_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__52_ccff_tail),
    .chany_top_out(sb_2__2__5_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__5_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__5_ccff_tail)
  );


  sb_2__2_
  sb_8__2_
  (
    .clk_2_N_in(clk_3_wires[43]),
    .clk_2_W_out(clk_2_wires[71]),
    .clk_2_E_out(clk_2_wires[69]),
    .prog_clk_2_N_in(prog_clk_3_wires[43]),
    .prog_clk_2_W_out(prog_clk_2_wires[71]),
    .prog_clk_2_E_out(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[299]),
    .config_enable_E_out(config_enableWires[143]),
    .config_enable_N_out(config_enableWires[142]),
    .config_enable_W_in(config_enableWires[140]),
    .pReset_E_out(pResetWires[143]),
    .pReset_N_out(pResetWires[142]),
    .pReset_W_in(pResetWires[140]),
    .chany_top_in(cby_2__3__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__73_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_81_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__71_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__64_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__64_ccff_tail),
    .chany_top_out(sb_2__2__6_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__6_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__6_ccff_tail)
  );


  sb_2__2_
  sb_8__9_
  (
    .clk_3_N_out(clk_3_wires[40]),
    .clk_3_S_in(clk_3_wires[37]),
    .prog_clk_3_N_out(prog_clk_3_wires[40]),
    .prog_clk_3_S_in(prog_clk_3_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[320]),
    .config_enable_E_out(config_enableWires[486]),
    .config_enable_N_out(config_enableWires[485]),
    .config_enable_W_in(config_enableWires[483]),
    .pReset_E_out(pResetWires[486]),
    .pReset_N_out(pResetWires[485]),
    .pReset_W_in(pResetWires[483]),
    .chany_top_in(cby_2__3__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__79_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_87_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__77_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__70_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__70_ccff_tail),
    .chany_top_out(sb_2__2__7_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__7_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__7_ccff_tail)
  );


  sb_2__2_
  sb_10__2_
  (
    .clk_2_N_in(clk_3_wires[87]),
    .clk_2_E_out(clk_2_wires[114]),
    .prog_clk_2_N_in(prog_clk_3_wires[87]),
    .prog_clk_2_E_out(prog_clk_2_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[375]),
    .config_enable_E_out(config_enableWires[151]),
    .config_enable_N_out(config_enableWires[150]),
    .config_enable_W_in(config_enableWires[148]),
    .pReset_E_out(pResetWires[151]),
    .pReset_N_out(pResetWires[150]),
    .pReset_W_in(pResetWires[148]),
    .chany_top_in(cby_2__3__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__91_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_101_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__91_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_91_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__82_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_91_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__82_ccff_tail),
    .chany_top_out(sb_2__2__8_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__8_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__8_ccff_tail)
  );


  sb_2__2_
  sb_10__9_
  (
    .clk_3_N_out(clk_3_wires[84]),
    .clk_3_S_in(clk_3_wires[81]),
    .prog_clk_3_N_out(prog_clk_3_wires[84]),
    .prog_clk_3_S_in(prog_clk_3_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[396]),
    .config_enable_E_out(config_enableWires[494]),
    .config_enable_N_out(config_enableWires[493]),
    .config_enable_W_in(config_enableWires[491]),
    .pReset_E_out(pResetWires[494]),
    .pReset_N_out(pResetWires[493]),
    .pReset_W_in(pResetWires[491]),
    .chany_top_in(cby_2__3__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .chanx_right_in(cbx_1__1__97_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_107_top_width_0_height_0_subtile_0__pin_O_5_upper),
    .chany_bottom_in(cby_1__1__97_chany_top_out[0:19]),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_97_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__88_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_97_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__88_ccff_tail),
    .chany_top_out(sb_2__2__9_chany_top_out[0:19]),
    .chanx_right_out(sb_2__2__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__2__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__2__9_chanx_left_out[0:19]),
    .ccff_tail(sb_2__2__9_ccff_tail)
  );


  sb_2__3_
  sb_2__3_
  (
    .clk_3_S_out(clk_3_wires[68]),
    .clk_3_N_in(clk_3_wires[65]),
    .prog_clk_3_S_out(prog_clk_3_wires[68]),
    .prog_clk_3_N_in(prog_clk_3_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[74]),
    .config_enable_E_in(config_enableWires[168]),
    .config_enable_N_out(config_enableWires[167]),
    .config_enable_W_out(config_enableWires[165]),
    .pReset_E_in(pResetWires[168]),
    .pReset_N_out(pResetWires[167]),
    .pReset_W_out(pResetWires[165]),
    .chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__2_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_2_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__0_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_0_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__0_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_0_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__0_ccff_tail),
    .chany_top_out(sb_2__3__0_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__0_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__0_ccff_tail)
  );


  sb_2__3_
  sb_2__10_
  (
    .clk_2_S_in(clk_3_wires[67]),
    .clk_2_W_out(clk_2_wires[21]),
    .prog_clk_2_S_in(prog_clk_3_wires[67]),
    .prog_clk_2_W_out(prog_clk_2_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[95]),
    .config_enable_E_in(config_enableWires[511]),
    .config_enable_N_out(config_enableWires[510]),
    .config_enable_W_out(config_enableWires[508]),
    .pReset_E_in(pResetWires[511]),
    .pReset_N_out(pResetWires[510]),
    .pReset_W_out(pResetWires[508]),
    .chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__3_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_3_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__1_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_1_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__1_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_1_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__1_ccff_tail),
    .chany_top_out(sb_2__3__1_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__1_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__1_ccff_tail)
  );


  sb_2__3_
  sb_4__3_
  (
    .clk_3_S_out(clk_3_wires[24]),
    .clk_3_N_in(clk_3_wires[21]),
    .prog_clk_3_S_out(prog_clk_3_wires[24]),
    .prog_clk_3_N_in(prog_clk_3_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[150]),
    .config_enable_E_in(config_enableWires[176]),
    .config_enable_N_out(config_enableWires[175]),
    .config_enable_W_out(config_enableWires[173]),
    .pReset_E_in(pResetWires[176]),
    .pReset_N_out(pResetWires[175]),
    .pReset_W_out(pResetWires[173]),
    .chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__4_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_4_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__2_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_2_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__2_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_2_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__2_ccff_tail),
    .chany_top_out(sb_2__3__2_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__2_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__2_ccff_tail)
  );


  sb_2__3_
  sb_4__10_
  (
    .clk_2_S_in(clk_3_wires[23]),
    .clk_2_W_out(clk_2_wires[62]),
    .clk_2_E_out(clk_2_wires[60]),
    .prog_clk_2_S_in(prog_clk_3_wires[23]),
    .prog_clk_2_W_out(prog_clk_2_wires[62]),
    .prog_clk_2_E_out(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[171]),
    .config_enable_E_in(config_enableWires[519]),
    .config_enable_N_out(config_enableWires[518]),
    .config_enable_W_out(config_enableWires[516]),
    .pReset_E_in(pResetWires[519]),
    .pReset_N_out(pResetWires[518]),
    .pReset_W_out(pResetWires[516]),
    .chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__5_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_5_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__3_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_3_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__3_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_3_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__3_ccff_tail),
    .chany_top_out(sb_2__3__3_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__3_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__3_ccff_tail)
  );


  sb_2__3_
  sb_6__3_
  (
    .clk_3_N_out(clk_3_wires[96]),
    .clk_3_S_in(clk_3_wires[93]),
    .prog_clk_3_N_out(prog_clk_3_wires[96]),
    .prog_clk_3_S_in(prog_clk_3_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[226]),
    .config_enable_E_out(config_enableWires[184]),
    .config_enable_W_out(config_enableWires[181]),
    .config_enable_N_out(config_enableWires[183]),
    .config_enable_S_in(config_enableWires[6]),
    .reset_N_out(resetWires[7]),
    .reset_S_in(resetWires[6]),
    .Test_en_N_out(Test_enWires[7]),
    .Test_en_S_in(Test_enWires[6]),
    .pReset_E_out(pResetWires[184]),
    .pReset_W_out(pResetWires[181]),
    .pReset_N_out(pResetWires[183]),
    .pReset_S_in(pResetWires[6]),
    .chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__6_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_6_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__4_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_4_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__4_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_4_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__4_ccff_tail),
    .chany_top_out(sb_2__3__4_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__4_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__4_ccff_tail)
  );


  sb_2__3_
  sb_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[247]),
    .config_enable_E_out(config_enableWires[527]),
    .config_enable_W_out(config_enableWires[524]),
    .config_enable_N_out(config_enableWires[526]),
    .config_enable_S_in(config_enableWires[20]),
    .reset_N_out(resetWires[21]),
    .reset_S_in(resetWires[20]),
    .Test_en_N_out(Test_enWires[21]),
    .Test_en_S_in(Test_enWires[20]),
    .pReset_E_out(pResetWires[527]),
    .pReset_W_out(pResetWires[524]),
    .pReset_N_out(pResetWires[526]),
    .pReset_S_in(pResetWires[20]),
    .chany_top_in(cby_1__1__58_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__7_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_7_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__5_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_5_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__5_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_5_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__5_ccff_tail),
    .chany_top_out(sb_2__3__5_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__5_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__5_ccff_tail)
  );


  sb_2__3_
  sb_8__3_
  (
    .clk_3_S_out(clk_3_wires[42]),
    .clk_3_N_in(clk_3_wires[39]),
    .prog_clk_3_S_out(prog_clk_3_wires[42]),
    .prog_clk_3_N_in(prog_clk_3_wires[39]),
    .prog_clk_0_N_in(prog_clk_0_wires[302]),
    .config_enable_E_out(config_enableWires[192]),
    .config_enable_N_out(config_enableWires[191]),
    .config_enable_W_in(config_enableWires[189]),
    .pReset_E_out(pResetWires[192]),
    .pReset_N_out(pResetWires[191]),
    .pReset_W_in(pResetWires[189]),
    .chany_top_in(cby_1__1__72_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__8_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_8_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__6_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_6_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__6_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_6_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__6_ccff_tail),
    .chany_top_out(sb_2__3__6_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__6_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__6_ccff_tail)
  );


  sb_2__3_
  sb_8__10_
  (
    .clk_2_S_in(clk_3_wires[41]),
    .clk_2_W_out(clk_2_wires[106]),
    .clk_2_E_out(clk_2_wires[104]),
    .prog_clk_2_S_in(prog_clk_3_wires[41]),
    .prog_clk_2_W_out(prog_clk_2_wires[106]),
    .prog_clk_2_E_out(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[323]),
    .config_enable_E_out(config_enableWires[535]),
    .config_enable_N_out(config_enableWires[534]),
    .config_enable_W_in(config_enableWires[532]),
    .pReset_E_out(pResetWires[535]),
    .pReset_N_out(pResetWires[534]),
    .pReset_W_in(pResetWires[532]),
    .chany_top_in(cby_1__1__78_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__9_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_9_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__7_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_7_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__7_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_7_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__7_ccff_tail),
    .chany_top_out(sb_2__3__7_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__7_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__7_ccff_tail)
  );


  sb_2__3_
  sb_10__3_
  (
    .clk_3_S_out(clk_3_wires[86]),
    .clk_3_N_in(clk_3_wires[83]),
    .prog_clk_3_S_out(prog_clk_3_wires[86]),
    .prog_clk_3_N_in(prog_clk_3_wires[83]),
    .prog_clk_0_N_in(prog_clk_0_wires[378]),
    .config_enable_E_out(config_enableWires[200]),
    .config_enable_N_out(config_enableWires[199]),
    .config_enable_W_in(config_enableWires[197]),
    .pReset_E_out(pResetWires[200]),
    .pReset_N_out(pResetWires[199]),
    .pReset_W_in(pResetWires[197]),
    .chany_top_in(cby_1__1__92_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_92_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__10_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_10_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__8_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_8_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__8_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_8_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__8_ccff_tail),
    .chany_top_out(sb_2__3__8_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__8_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__8_ccff_tail)
  );


  sb_2__3_
  sb_10__10_
  (
    .clk_2_S_in(clk_3_wires[85]),
    .clk_2_E_out(clk_2_wires[133]),
    .prog_clk_2_S_in(prog_clk_3_wires[85]),
    .prog_clk_2_E_out(prog_clk_2_wires[133]),
    .prog_clk_0_N_in(prog_clk_0_wires[399]),
    .config_enable_E_out(config_enableWires[543]),
    .config_enable_N_out(config_enableWires[542]),
    .config_enable_W_in(config_enableWires[540]),
    .pReset_E_out(pResetWires[543]),
    .pReset_N_out(pResetWires[542]),
    .pReset_W_in(pResetWires[540]),
    .chany_top_in(cby_1__1__98_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_98_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .chanx_right_in(cbx_1__3__11_chanx_left_out[0:19]),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_0_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_1_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_2_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_3_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_4_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_5_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_6_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_7_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_8_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_9_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_10_upper),
    .right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_11_top_width_0_height_0_subtile_0__pin_out_11_upper),
    .chany_bottom_in(cby_2__3__9_chany_top_out[0:19]),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_9_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__9_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_9_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__9_ccff_tail),
    .chany_top_out(sb_2__3__9_chany_top_out[0:19]),
    .chanx_right_out(sb_2__3__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_2__3__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_2__3__9_chanx_left_out[0:19]),
    .ccff_tail(sb_2__3__9_ccff_tail)
  );


  sb_4__0_
  sb_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[445]),
    .config_enable_N_out(config_enableWires[60]),
    .config_enable_W_in(config_enableWires[59]),
    .pReset_N_out(pResetWires[60]),
    .pReset_W_in(pResetWires[59]),
    .chany_top_in(cby_12__1__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chanx_left_in(cbx_1__0__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_head(grid_io_bottom_bottom_0_ccff_tail),
    .chany_top_out(sb_12__0__0_chany_top_out[0:19]),
    .chanx_left_out(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[11])
  );


  sb_4__1_
  sb_12__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[448]),
    .config_enable_N_out(config_enableWires[109]),
    .config_enable_W_in(config_enableWires[107]),
    .pReset_N_out(pResetWires[109]),
    .pReset_W_in(pResetWires[107]),
    .chany_top_in(cby_12__1__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__0_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_110_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__99_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_110_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__99_ccff_tail),
    .chany_top_out(sb_12__1__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[10])
  );


  sb_4__1_
  sb_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[457]),
    .config_enable_N_out(config_enableWires[256]),
    .config_enable_W_in(config_enableWires[254]),
    .pReset_N_out(pResetWires[256]),
    .pReset_W_in(pResetWires[254]),
    .chany_top_in(cby_12__1__3_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__2_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__101_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_112_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__101_ccff_tail),
    .chany_top_out(sb_12__1__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[7])
  );


  sb_4__1_
  sb_12__5_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[460]),
    .config_enable_N_out(config_enableWires[305]),
    .config_enable_W_in(config_enableWires[303]),
    .pReset_N_out(pResetWires[305]),
    .pReset_W_in(pResetWires[303]),
    .chany_top_in(cby_12__1__4_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__3_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_113_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__102_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_113_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__102_ccff_tail),
    .chany_top_out(sb_12__1__2_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[6])
  );


  sb_4__1_
  sb_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[463]),
    .config_enable_N_out(config_enableWires[354]),
    .config_enable_W_in(config_enableWires[352]),
    .pReset_N_out(pResetWires[354]),
    .pReset_W_in(pResetWires[352]),
    .chany_top_in(cby_12__1__5_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__4_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_114_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__103_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_114_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__103_ccff_tail),
    .chany_top_out(sb_12__1__3_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[5])
  );


  sb_4__1_
  sb_12__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[466]),
    .config_enable_N_out(config_enableWires[403]),
    .config_enable_W_in(config_enableWires[401]),
    .pReset_N_out(pResetWires[403]),
    .pReset_W_in(pResetWires[401]),
    .chany_top_in(cby_12__1__6_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__5_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_115_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__104_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_115_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__104_ccff_tail),
    .chany_top_out(sb_12__1__4_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[4])
  );


  sb_4__1_
  sb_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[469]),
    .config_enable_N_out(config_enableWires[452]),
    .config_enable_W_in(config_enableWires[450]),
    .pReset_N_out(pResetWires[452]),
    .pReset_W_in(pResetWires[450]),
    .chany_top_in(cby_12__1__7_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__6_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_116_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__105_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_116_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__105_ccff_tail),
    .chany_top_out(sb_12__1__5_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[3])
  );


  sb_4__1_
  sb_12__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[478]),
    .config_enable_N_out(config_enableWires[599]),
    .config_enable_W_in(config_enableWires[597]),
    .pReset_N_out(pResetWires[599]),
    .pReset_W_in(pResetWires[597]),
    .chany_top_in(cby_12__1__9_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__8_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__107_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_118_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__107_ccff_tail),
    .chany_top_out(sb_12__1__6_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[0])
  );


  sb_4__2_
  sb_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[451]),
    .config_enable_N_out(config_enableWires[158]),
    .config_enable_W_in(config_enableWires[156]),
    .pReset_N_out(pResetWires[158]),
    .pReset_W_in(pResetWires[156]),
    .chany_top_in(cby_12__3__0_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__1_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_111_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__100_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_111_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__100_ccff_tail),
    .chany_top_out(sb_12__2__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__2__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__2__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[9])
  );


  sb_4__2_
  sb_12__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[472]),
    .config_enable_N_out(config_enableWires[501]),
    .config_enable_W_in(config_enableWires[499]),
    .pReset_N_out(pResetWires[501]),
    .pReset_W_in(pResetWires[499]),
    .chany_top_in(cby_12__3__1_chany_bottom_out[0:19]),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_lower),
    .top_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__1__7_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_117_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__1__106_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_117_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(cbx_1__1__106_ccff_tail),
    .chany_top_out(sb_12__2__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__2__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__2__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[2])
  );


  sb_4__3_
  sb_12__3_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[454]),
    .config_enable_N_out(config_enableWires[207]),
    .config_enable_W_in(config_enableWires[205]),
    .pReset_N_out(pResetWires[207]),
    .pReset_W_in(pResetWires[205]),
    .chany_top_in(cby_12__1__2_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_112_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__3__0_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_10_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__10_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_10_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__10_ccff_tail),
    .chany_top_out(sb_12__3__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__3__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__3__0_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[8])
  );


  sb_4__3_
  sb_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[475]),
    .config_enable_N_out(config_enableWires[550]),
    .config_enable_W_in(config_enableWires[548]),
    .pReset_N_out(pResetWires[550]),
    .pReset_W_in(pResetWires[548]),
    .chany_top_in(cby_12__1__8_chany_bottom_out[0:19]),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_6_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_7_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_8_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_9_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_10_lower),
    .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_118_right_width_0_height_0_subtile_0__pin_O_11_lower),
    .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .chany_bottom_in(cby_12__3__1_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_24_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_24_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_25_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_25_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_26_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_26_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_27_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_27_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_28_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_28_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_29_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_29_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_30_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_30_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_31_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_31_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_32_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_32_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_33_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_33_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_34_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_34_upper),
    .bottom_left_grid_right_width_1_height_0_subtile_0__pin_out_35_(grid_mult_18_11_right_width_1_height_0_subtile_0__pin_out_35_upper),
    .chanx_left_in(cbx_2__3__11_chanx_right_out[0:19]),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_12_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_12_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_13_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_13_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_14_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_14_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_15_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_15_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_16_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_16_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_17_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_17_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_18_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_18_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_19_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_19_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_20_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_20_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_21_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_21_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_22_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_22_lower),
    .left_bottom_grid_top_width_1_height_0_subtile_0__pin_out_23_(grid_mult_18_11_top_width_1_height_0_subtile_0__pin_out_23_lower),
    .ccff_head(cbx_2__3__11_ccff_tail),
    .chany_top_out(sb_12__3__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__3__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__3__1_chanx_left_out[0:19]),
    .ccff_tail(ccff_tail[1])
  );


  sb_4__4_
  sb_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[480]),
    .sc_head_E_out(sc_tail),
    .config_enable_W_in(config_enableWires[635]),
    .sc_head_W_in(sc_headWires[312]),
    .pReset_W_in(pResetWires[635]),
    .chany_bottom_in(cby_12__1__9_chany_top_out[0:19]),
    .bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_6_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_7_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_8_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_9_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_10_upper),
    .bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_119_right_width_0_height_0_subtile_0__pin_O_11_upper),
    .chanx_left_in(cbx_1__12__11_chanx_right_out[0:19]),
    .left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_0_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_1_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_2_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_3_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_4_lower),
    .left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_119_top_width_0_height_0_subtile_0__pin_O_5_lower),
    .ccff_head(ccff_head[0]),
    .chany_bottom_out(sb_12__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_12__12__0_ccff_tail)
  );


  cbx_1__0_
  cbx_1__0_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[0]),
    .config_enable_E_in(config_enableWires[26]),
    .config_enable_W_out(config_enableWires[25]),
    .sc_head_E_out(sc_headWires[26]),
    .sc_head_N_in(sc_headWires[25]),
    .pReset_E_in(pResetWires[26]),
    .pReset_W_out(pResetWires[25]),
    .chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__0__0_ccff_tail),
    .chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[123:131]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[123:131]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[123:131]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_11_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_11_ccff_tail)
  );


  cbx_1__0_
  cbx_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[63]),
    .config_enable_E_in(config_enableWires[29]),
    .config_enable_W_out(config_enableWires[28]),
    .sc_head_N_out(sc_headWires[28]),
    .sc_head_W_in(sc_headWires[27]),
    .pReset_E_in(pResetWires[29]),
    .pReset_W_out(pResetWires[28]),
    .chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__0_ccff_tail),
    .chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[114:122]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[114:122]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[114:122]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_10_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_10_ccff_tail)
  );


  cbx_1__0_
  cbx_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[101]),
    .config_enable_E_in(config_enableWires[32]),
    .config_enable_W_out(config_enableWires[31]),
    .sc_head_E_out(sc_headWires[78]),
    .sc_head_N_in(sc_headWires[77]),
    .pReset_E_in(pResetWires[32]),
    .pReset_W_out(pResetWires[31]),
    .chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__1_ccff_tail),
    .chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[105:113]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[105:113]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[105:113]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_9_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_9_ccff_tail)
  );


  cbx_1__0_
  cbx_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[139]),
    .config_enable_E_in(config_enableWires[35]),
    .config_enable_W_out(config_enableWires[34]),
    .sc_head_N_out(sc_headWires[80]),
    .sc_head_W_in(sc_headWires[79]),
    .pReset_E_in(pResetWires[35]),
    .pReset_W_out(pResetWires[34]),
    .chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__2_ccff_tail),
    .chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[96:104]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[96:104]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[96:104]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_8_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_8_ccff_tail)
  );


  cbx_1__0_
  cbx_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[177]),
    .config_enable_E_in(config_enableWires[38]),
    .config_enable_W_out(config_enableWires[37]),
    .sc_head_E_out(sc_headWires[130]),
    .sc_head_N_in(sc_headWires[129]),
    .pReset_E_in(pResetWires[38]),
    .pReset_W_out(pResetWires[37]),
    .chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__3_ccff_tail),
    .chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[87:95]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[87:95]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[87:95]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_7_ccff_tail)
  );


  cbx_1__0_
  cbx_6__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[215]),
    .config_enable_E_in(config_enableWires[41]),
    .config_enable_W_out(config_enableWires[40]),
    .sc_head_N_out(sc_headWires[132]),
    .sc_head_W_in(sc_headWires[131]),
    .pReset_E_in(pResetWires[41]),
    .pReset_W_out(pResetWires[40]),
    .chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__4_ccff_tail),
    .chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[78:86]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[78:86]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[78:86]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_6_ccff_tail)
  );


  cbx_1__0_
  cbx_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[253]),
    .config_enable_E_out(config_enableWires[44]),
    .config_enable_W_in(config_enableWires[43]),
    .sc_head_E_out(sc_headWires[182]),
    .sc_head_N_in(sc_headWires[181]),
    .pReset_E_out(pResetWires[44]),
    .pReset_W_in(pResetWires[43]),
    .chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__5_ccff_tail),
    .chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[69:77]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[69:77]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[69:77]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_5_ccff_tail)
  );


  cbx_1__0_
  cbx_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[291]),
    .config_enable_E_out(config_enableWires[47]),
    .config_enable_W_in(config_enableWires[46]),
    .sc_head_N_out(sc_headWires[184]),
    .sc_head_W_in(sc_headWires[183]),
    .pReset_E_out(pResetWires[47]),
    .pReset_W_in(pResetWires[46]),
    .chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__6_ccff_tail),
    .chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[60:68]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[60:68]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[60:68]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_4_ccff_tail)
  );


  cbx_1__0_
  cbx_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[329]),
    .config_enable_E_out(config_enableWires[50]),
    .config_enable_W_in(config_enableWires[49]),
    .sc_head_E_out(sc_headWires[234]),
    .sc_head_N_in(sc_headWires[233]),
    .pReset_E_out(pResetWires[50]),
    .pReset_W_in(pResetWires[49]),
    .chanx_left_in(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__7_ccff_tail),
    .chanx_left_out(cbx_1__0__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__8_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[51:59]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[51:59]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[51:59]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_3_ccff_tail)
  );


  cbx_1__0_
  cbx_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[367]),
    .config_enable_E_out(config_enableWires[53]),
    .config_enable_W_in(config_enableWires[52]),
    .sc_head_N_out(sc_headWires[236]),
    .sc_head_W_in(sc_headWires[235]),
    .pReset_E_out(pResetWires[53]),
    .pReset_W_in(pResetWires[52]),
    .chanx_left_in(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__8_ccff_tail),
    .chanx_left_out(cbx_1__0__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__9_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[42:50]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[42:50]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[42:50]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_2_ccff_tail)
  );


  cbx_1__0_
  cbx_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[405]),
    .config_enable_E_out(config_enableWires[56]),
    .config_enable_W_in(config_enableWires[55]),
    .sc_head_E_out(sc_headWires[286]),
    .sc_head_N_in(sc_headWires[285]),
    .pReset_E_out(pResetWires[56]),
    .pReset_W_in(pResetWires[55]),
    .chanx_left_in(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__9_ccff_tail),
    .chanx_left_out(cbx_1__0__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__10_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[33:41]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[33:41]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[33:41]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_1_ccff_tail)
  );


  cbx_1__0_
  cbx_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[443]),
    .config_enable_E_out(config_enableWires[59]),
    .config_enable_W_in(config_enableWires[58]),
    .sc_head_N_out(sc_headWires[288]),
    .sc_head_W_in(sc_headWires[287]),
    .pReset_E_out(pResetWires[59]),
    .pReset_W_in(pResetWires[58]),
    .chanx_left_in(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__10_ccff_tail),
    .chanx_left_out(cbx_1__0__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__11_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[24:32]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[24:32]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[24:32]),
    .top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
    .top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
    .top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
    .ccff_tail(grid_io_bottom_bottom_0_ccff_tail)
  );


  cbx_1__1_
  cbx_1__1_
  (
    .clk_1_S_out(clk_1_wires[4]),
    .clk_1_N_out(clk_1_wires[3]),
    .clk_1_E_in(clk_1_wires[2]),
    .prog_clk_1_S_out(prog_clk_1_wires[4]),
    .prog_clk_1_N_out(prog_clk_1_wires[3]),
    .prog_clk_1_E_in(prog_clk_1_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[6]),
    .prog_clk_0_W_out(prog_clk_0_wires[4]),
    .config_enable_S_out(config_enableWires[63]),
    .config_enable_E_in(config_enableWires[62]),
    .config_enable_W_out(config_enableWires[61]),
    .sc_head_S_out(sc_headWires[24]),
    .sc_head_N_in(sc_headWires[23]),
    .pReset_S_out(pResetWires[63]),
    .pReset_E_in(pResetWires[62]),
    .pReset_W_out(pResetWires[61]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[0]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[0]),
    .chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__0_ccff_tail),
    .chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__0_ccff_tail)
  );


  cbx_1__1_
  cbx_1__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[10]),
    .config_enable_S_out(config_enableWires[112]),
    .config_enable_E_in(config_enableWires[111]),
    .config_enable_W_out(config_enableWires[110]),
    .sc_head_S_out(sc_headWires[22]),
    .sc_head_N_in(sc_headWires[21]),
    .pReset_S_out(pResetWires[112]),
    .pReset_E_in(pResetWires[111]),
    .pReset_W_out(pResetWires[110]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[1]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[1]),
    .chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__1_ccff_tail),
    .chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__1_ccff_tail)
  );


  cbx_1__1_
  cbx_1__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[21]),
    .prog_clk_0_W_out(prog_clk_0_wires[20]),
    .config_enable_S_out(config_enableWires[210]),
    .config_enable_E_in(config_enableWires[209]),
    .config_enable_W_out(config_enableWires[208]),
    .sc_head_S_out(sc_headWires[18]),
    .sc_head_N_in(sc_headWires[17]),
    .pReset_S_out(pResetWires[210]),
    .pReset_E_in(pResetWires[209]),
    .pReset_W_out(pResetWires[208]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[3]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[3]),
    .chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__2_ccff_tail),
    .chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__2_ccff_tail)
  );


  cbx_1__1_
  cbx_1__5_
  (
    .clk_1_S_out(clk_1_wires[18]),
    .clk_1_N_out(clk_1_wires[17]),
    .clk_1_E_in(clk_1_wires[16]),
    .prog_clk_1_S_out(prog_clk_1_wires[18]),
    .prog_clk_1_N_out(prog_clk_1_wires[17]),
    .prog_clk_1_E_in(prog_clk_1_wires[16]),
    .prog_clk_0_N_in(prog_clk_0_wires[26]),
    .prog_clk_0_W_out(prog_clk_0_wires[25]),
    .config_enable_S_out(config_enableWires[259]),
    .config_enable_E_in(config_enableWires[258]),
    .config_enable_W_out(config_enableWires[257]),
    .sc_head_S_out(sc_headWires[16]),
    .sc_head_N_in(sc_headWires[15]),
    .pReset_S_out(pResetWires[259]),
    .pReset_E_in(pResetWires[258]),
    .pReset_W_out(pResetWires[257]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[4]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[4]),
    .chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__3_ccff_tail),
    .chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__3_ccff_tail)
  );


  cbx_1__1_
  cbx_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[30]),
    .config_enable_S_out(config_enableWires[308]),
    .config_enable_E_in(config_enableWires[307]),
    .config_enable_W_out(config_enableWires[306]),
    .sc_head_S_out(sc_headWires[14]),
    .sc_head_N_in(sc_headWires[13]),
    .pReset_S_out(pResetWires[308]),
    .pReset_E_in(pResetWires[307]),
    .pReset_W_out(pResetWires[306]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[5]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[5]),
    .chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__4_ccff_tail),
    .chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__4_ccff_tail)
  );


  cbx_1__1_
  cbx_1__7_
  (
    .clk_1_S_out(clk_1_wires[25]),
    .clk_1_N_out(clk_1_wires[24]),
    .clk_1_E_in(clk_1_wires[23]),
    .prog_clk_1_S_out(prog_clk_1_wires[25]),
    .prog_clk_1_N_out(prog_clk_1_wires[24]),
    .prog_clk_1_E_in(prog_clk_1_wires[23]),
    .prog_clk_0_N_in(prog_clk_0_wires[36]),
    .prog_clk_0_W_out(prog_clk_0_wires[35]),
    .config_enable_S_out(config_enableWires[357]),
    .config_enable_E_in(config_enableWires[356]),
    .config_enable_W_out(config_enableWires[355]),
    .sc_head_S_out(sc_headWires[12]),
    .sc_head_N_in(sc_headWires[11]),
    .pReset_S_out(pResetWires[357]),
    .pReset_E_in(pResetWires[356]),
    .pReset_W_out(pResetWires[355]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[6]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[6]),
    .chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__5_ccff_tail),
    .chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__5_ccff_tail)
  );


  cbx_1__1_
  cbx_1__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[41]),
    .prog_clk_0_W_out(prog_clk_0_wires[40]),
    .config_enable_S_out(config_enableWires[406]),
    .config_enable_E_in(config_enableWires[405]),
    .config_enable_W_out(config_enableWires[404]),
    .sc_head_S_out(sc_headWires[10]),
    .sc_head_N_in(sc_headWires[9]),
    .pReset_S_out(pResetWires[406]),
    .pReset_E_in(pResetWires[405]),
    .pReset_W_out(pResetWires[404]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[7]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[7]),
    .chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__6_ccff_tail),
    .chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__6_ccff_tail)
  );


  cbx_1__1_
  cbx_1__9_
  (
    .clk_1_S_out(clk_1_wires[32]),
    .clk_1_N_out(clk_1_wires[31]),
    .clk_1_E_in(clk_1_wires[30]),
    .prog_clk_1_S_out(prog_clk_1_wires[32]),
    .prog_clk_1_N_out(prog_clk_1_wires[31]),
    .prog_clk_1_E_in(prog_clk_1_wires[30]),
    .prog_clk_0_N_in(prog_clk_0_wires[46]),
    .prog_clk_0_W_out(prog_clk_0_wires[45]),
    .config_enable_S_out(config_enableWires[455]),
    .config_enable_E_in(config_enableWires[454]),
    .config_enable_W_out(config_enableWires[453]),
    .sc_head_S_out(sc_headWires[8]),
    .sc_head_N_in(sc_headWires[7]),
    .pReset_S_out(pResetWires[455]),
    .pReset_E_in(pResetWires[454]),
    .pReset_W_out(pResetWires[453]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[8]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[8]),
    .chanx_left_in(sb_0__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__7_ccff_tail),
    .chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__7_ccff_tail)
  );


  cbx_1__1_
  cbx_1__11_
  (
    .clk_1_S_out(clk_1_wires[39]),
    .clk_1_N_out(clk_1_wires[38]),
    .clk_1_E_in(clk_1_wires[37]),
    .prog_clk_1_S_out(prog_clk_1_wires[39]),
    .prog_clk_1_N_out(prog_clk_1_wires[38]),
    .prog_clk_1_E_in(prog_clk_1_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[56]),
    .prog_clk_0_W_out(prog_clk_0_wires[55]),
    .config_enable_S_out(config_enableWires[553]),
    .config_enable_E_in(config_enableWires[552]),
    .config_enable_W_out(config_enableWires[551]),
    .sc_head_S_out(sc_headWires[4]),
    .sc_head_N_in(sc_headWires[3]),
    .pReset_S_out(pResetWires[553]),
    .pReset_E_in(pResetWires[552]),
    .pReset_W_out(pResetWires[551]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[10]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[10]),
    .chanx_left_in(sb_0__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_0__1__8_ccff_tail),
    .chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__8_ccff_tail)
  );


  cbx_1__1_
  cbx_2__1_
  (
    .clk_1_S_out(clk_1_wires[6]),
    .clk_1_N_out(clk_1_wires[5]),
    .clk_1_W_in(clk_1_wires[1]),
    .prog_clk_1_S_out(prog_clk_1_wires[6]),
    .prog_clk_1_N_out(prog_clk_1_wires[5]),
    .prog_clk_1_W_in(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[66]),
    .config_enable_S_out(config_enableWires[68]),
    .config_enable_E_in(config_enableWires[67]),
    .config_enable_W_out(config_enableWires[66]),
    .sc_head_N_out(sc_headWires[30]),
    .sc_head_S_in(sc_headWires[29]),
    .pReset_S_out(pResetWires[68]),
    .pReset_E_in(pResetWires[67]),
    .pReset_W_out(pResetWires[66]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[11]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[11]),
    .chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__0_ccff_tail),
    .chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__9_ccff_tail)
  );


  cbx_1__1_
  cbx_2__2_
  (
    .clk_2_E_in(clk_2_wires[2]),
    .clk_2_W_out(clk_2_wires[1]),
    .prog_clk_2_E_in(prog_clk_2_wires[2]),
    .prog_clk_2_W_out(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[69]),
    .config_enable_S_out(config_enableWires[117]),
    .config_enable_E_in(config_enableWires[116]),
    .config_enable_W_out(config_enableWires[115]),
    .sc_head_N_out(sc_headWires[32]),
    .sc_head_S_in(sc_headWires[31]),
    .pReset_S_out(pResetWires[117]),
    .pReset_E_in(pResetWires[116]),
    .pReset_W_out(pResetWires[115]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[12]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[12]),
    .chanx_left_in(sb_1__2__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__0_ccff_tail),
    .chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__10_ccff_tail)
  );


  cbx_1__1_
  cbx_2__4_
  (
    .clk_2_E_in(clk_2_wires[7]),
    .clk_2_W_out(clk_2_wires[6]),
    .prog_clk_2_E_in(prog_clk_2_wires[7]),
    .prog_clk_2_W_out(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[75]),
    .config_enable_S_out(config_enableWires[215]),
    .config_enable_E_in(config_enableWires[214]),
    .config_enable_W_out(config_enableWires[213]),
    .sc_head_N_out(sc_headWires[36]),
    .sc_head_S_in(sc_headWires[35]),
    .pReset_S_out(pResetWires[215]),
    .pReset_E_in(pResetWires[214]),
    .pReset_W_out(pResetWires[213]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[14]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[14]),
    .chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__1_ccff_tail),
    .chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__11_ccff_tail)
  );


  cbx_1__1_
  cbx_2__5_
  (
    .clk_1_S_out(clk_1_wires[20]),
    .clk_1_N_out(clk_1_wires[19]),
    .clk_1_W_in(clk_1_wires[15]),
    .prog_clk_1_S_out(prog_clk_1_wires[20]),
    .prog_clk_1_N_out(prog_clk_1_wires[19]),
    .prog_clk_1_W_in(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[78]),
    .config_enable_S_out(config_enableWires[264]),
    .config_enable_E_in(config_enableWires[263]),
    .config_enable_W_out(config_enableWires[262]),
    .sc_head_N_out(sc_headWires[38]),
    .sc_head_S_in(sc_headWires[37]),
    .pReset_S_out(pResetWires[264]),
    .pReset_E_in(pResetWires[263]),
    .pReset_W_out(pResetWires[262]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[15]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[15]),
    .chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__2_ccff_tail),
    .chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__12_ccff_tail)
  );


  cbx_1__1_
  cbx_2__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[81]),
    .config_enable_S_out(config_enableWires[313]),
    .config_enable_E_in(config_enableWires[312]),
    .config_enable_W_out(config_enableWires[311]),
    .sc_head_N_out(sc_headWires[40]),
    .sc_head_S_in(sc_headWires[39]),
    .pReset_S_out(pResetWires[313]),
    .pReset_E_in(pResetWires[312]),
    .pReset_W_out(pResetWires[311]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[16]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[16]),
    .chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__3_ccff_tail),
    .chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__13_ccff_tail)
  );


  cbx_1__1_
  cbx_2__7_
  (
    .clk_1_S_out(clk_1_wires[27]),
    .clk_1_N_out(clk_1_wires[26]),
    .clk_1_W_in(clk_1_wires[22]),
    .prog_clk_1_S_out(prog_clk_1_wires[27]),
    .prog_clk_1_N_out(prog_clk_1_wires[26]),
    .prog_clk_1_W_in(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[84]),
    .config_enable_S_out(config_enableWires[362]),
    .config_enable_E_in(config_enableWires[361]),
    .config_enable_W_out(config_enableWires[360]),
    .sc_head_N_out(sc_headWires[42]),
    .sc_head_S_in(sc_headWires[41]),
    .pReset_S_out(pResetWires[362]),
    .pReset_E_in(pResetWires[361]),
    .pReset_W_out(pResetWires[360]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[17]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[17]),
    .chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__4_ccff_tail),
    .chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__14_ccff_tail)
  );


  cbx_1__1_
  cbx_2__8_
  (
    .clk_2_E_in(clk_2_wires[14]),
    .clk_2_W_out(clk_2_wires[13]),
    .prog_clk_2_E_in(prog_clk_2_wires[14]),
    .prog_clk_2_W_out(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[87]),
    .config_enable_S_out(config_enableWires[411]),
    .config_enable_E_in(config_enableWires[410]),
    .config_enable_W_out(config_enableWires[409]),
    .sc_head_N_out(sc_headWires[44]),
    .sc_head_S_in(sc_headWires[43]),
    .pReset_S_out(pResetWires[411]),
    .pReset_E_in(pResetWires[410]),
    .pReset_W_out(pResetWires[409]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[18]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[18]),
    .chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__5_ccff_tail),
    .chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__15_ccff_tail)
  );


  cbx_1__1_
  cbx_2__9_
  (
    .clk_1_S_out(clk_1_wires[34]),
    .clk_1_N_out(clk_1_wires[33]),
    .clk_1_W_in(clk_1_wires[29]),
    .prog_clk_1_S_out(prog_clk_1_wires[34]),
    .prog_clk_1_N_out(prog_clk_1_wires[33]),
    .prog_clk_1_W_in(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[90]),
    .config_enable_S_out(config_enableWires[460]),
    .config_enable_E_in(config_enableWires[459]),
    .config_enable_W_out(config_enableWires[458]),
    .sc_head_N_out(sc_headWires[46]),
    .sc_head_S_in(sc_headWires[45]),
    .pReset_S_out(pResetWires[460]),
    .pReset_E_in(pResetWires[459]),
    .pReset_W_out(pResetWires[458]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[19]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[19]),
    .chanx_left_in(sb_1__2__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__1_ccff_tail),
    .chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__16_ccff_tail)
  );


  cbx_1__1_
  cbx_2__11_
  (
    .clk_1_S_out(clk_1_wires[41]),
    .clk_1_N_out(clk_1_wires[40]),
    .clk_1_W_in(clk_1_wires[36]),
    .prog_clk_1_S_out(prog_clk_1_wires[41]),
    .prog_clk_1_N_out(prog_clk_1_wires[40]),
    .prog_clk_1_W_in(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[96]),
    .config_enable_S_out(config_enableWires[558]),
    .config_enable_E_in(config_enableWires[557]),
    .config_enable_W_out(config_enableWires[556]),
    .sc_head_N_out(sc_headWires[50]),
    .sc_head_S_in(sc_headWires[49]),
    .pReset_S_out(pResetWires[558]),
    .pReset_E_in(pResetWires[557]),
    .pReset_W_out(pResetWires[556]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[21]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[21]),
    .chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__6_ccff_tail),
    .chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__17_ccff_tail)
  );


  cbx_1__1_
  cbx_3__1_
  (
    .clk_1_S_out(clk_1_wires[46]),
    .clk_1_N_out(clk_1_wires[45]),
    .clk_1_E_in(clk_1_wires[44]),
    .prog_clk_1_S_out(prog_clk_1_wires[46]),
    .prog_clk_1_N_out(prog_clk_1_wires[45]),
    .prog_clk_1_E_in(prog_clk_1_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[104]),
    .config_enable_S_out(config_enableWires[72]),
    .config_enable_E_in(config_enableWires[71]),
    .config_enable_W_out(config_enableWires[70]),
    .sc_head_S_out(sc_headWires[76]),
    .sc_head_N_in(sc_headWires[75]),
    .pReset_S_out(pResetWires[72]),
    .pReset_E_in(pResetWires[71]),
    .pReset_W_out(pResetWires[70]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[22]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[22]),
    .chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__7_ccff_tail),
    .chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__18_ccff_tail)
  );


  cbx_1__1_
  cbx_3__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[107]),
    .config_enable_S_out(config_enableWires[121]),
    .config_enable_E_in(config_enableWires[120]),
    .config_enable_W_out(config_enableWires[119]),
    .sc_head_S_out(sc_headWires[74]),
    .sc_head_N_in(sc_headWires[73]),
    .pReset_S_out(pResetWires[121]),
    .pReset_E_in(pResetWires[120]),
    .pReset_W_out(pResetWires[119]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[23]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[23]),
    .chanx_left_in(sb_2__2__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__2_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__0_ccff_tail),
    .chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__19_ccff_tail)
  );


  cbx_1__1_
  cbx_3__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[113]),
    .config_enable_S_out(config_enableWires[219]),
    .config_enable_E_in(config_enableWires[218]),
    .config_enable_W_out(config_enableWires[217]),
    .sc_head_S_out(sc_headWires[70]),
    .sc_head_N_in(sc_headWires[69]),
    .pReset_S_out(pResetWires[219]),
    .pReset_E_in(pResetWires[218]),
    .pReset_W_out(pResetWires[217]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[25]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[25]),
    .chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__8_ccff_tail),
    .chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__20_ccff_tail)
  );


  cbx_1__1_
  cbx_3__5_
  (
    .clk_1_S_out(clk_1_wires[60]),
    .clk_1_N_out(clk_1_wires[59]),
    .clk_1_E_in(clk_1_wires[58]),
    .prog_clk_1_S_out(prog_clk_1_wires[60]),
    .prog_clk_1_N_out(prog_clk_1_wires[59]),
    .prog_clk_1_E_in(prog_clk_1_wires[58]),
    .prog_clk_0_N_in(prog_clk_0_wires[116]),
    .config_enable_S_out(config_enableWires[268]),
    .config_enable_E_in(config_enableWires[267]),
    .config_enable_W_out(config_enableWires[266]),
    .sc_head_S_out(sc_headWires[68]),
    .sc_head_N_in(sc_headWires[67]),
    .pReset_S_out(pResetWires[268]),
    .pReset_E_in(pResetWires[267]),
    .pReset_W_out(pResetWires[266]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[26]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[26]),
    .chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__9_ccff_tail),
    .chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__21_ccff_tail)
  );


  cbx_1__1_
  cbx_3__6_
  (
    .clk_3_W_out(clk_3_wires[51]),
    .clk_3_E_in(clk_3_wires[50]),
    .prog_clk_3_W_out(prog_clk_3_wires[51]),
    .prog_clk_3_E_in(prog_clk_3_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[119]),
    .config_enable_S_out(config_enableWires[317]),
    .config_enable_E_in(config_enableWires[316]),
    .config_enable_W_out(config_enableWires[315]),
    .sc_head_S_out(sc_headWires[66]),
    .sc_head_N_in(sc_headWires[65]),
    .pReset_S_out(pResetWires[317]),
    .pReset_E_in(pResetWires[316]),
    .pReset_W_out(pResetWires[315]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[27]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[27]),
    .chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__10_ccff_tail),
    .chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__22_ccff_tail)
  );


  cbx_1__1_
  cbx_3__7_
  (
    .clk_1_S_out(clk_1_wires[67]),
    .clk_1_N_out(clk_1_wires[66]),
    .clk_1_E_in(clk_1_wires[65]),
    .prog_clk_1_S_out(prog_clk_1_wires[67]),
    .prog_clk_1_N_out(prog_clk_1_wires[66]),
    .prog_clk_1_E_in(prog_clk_1_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[122]),
    .config_enable_S_out(config_enableWires[366]),
    .config_enable_E_in(config_enableWires[365]),
    .config_enable_W_out(config_enableWires[364]),
    .sc_head_S_out(sc_headWires[64]),
    .sc_head_N_in(sc_headWires[63]),
    .pReset_S_out(pResetWires[366]),
    .pReset_E_in(pResetWires[365]),
    .pReset_W_out(pResetWires[364]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[28]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[28]),
    .chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__11_ccff_tail),
    .chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__23_ccff_tail)
  );


  cbx_1__1_
  cbx_3__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[125]),
    .config_enable_S_out(config_enableWires[415]),
    .config_enable_E_in(config_enableWires[414]),
    .config_enable_W_out(config_enableWires[413]),
    .sc_head_S_out(sc_headWires[62]),
    .sc_head_N_in(sc_headWires[61]),
    .pReset_S_out(pResetWires[415]),
    .pReset_E_in(pResetWires[414]),
    .pReset_W_out(pResetWires[413]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[29]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[29]),
    .chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__12_ccff_tail),
    .chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__24_ccff_tail)
  );


  cbx_1__1_
  cbx_3__9_
  (
    .clk_1_S_out(clk_1_wires[74]),
    .clk_1_N_out(clk_1_wires[73]),
    .clk_1_E_in(clk_1_wires[72]),
    .prog_clk_1_S_out(prog_clk_1_wires[74]),
    .prog_clk_1_N_out(prog_clk_1_wires[73]),
    .prog_clk_1_E_in(prog_clk_1_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[128]),
    .config_enable_S_out(config_enableWires[464]),
    .config_enable_E_in(config_enableWires[463]),
    .config_enable_W_out(config_enableWires[462]),
    .sc_head_S_out(sc_headWires[60]),
    .sc_head_N_in(sc_headWires[59]),
    .pReset_S_out(pResetWires[464]),
    .pReset_E_in(pResetWires[463]),
    .pReset_W_out(pResetWires[462]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[30]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[30]),
    .chanx_left_in(sb_2__2__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__3_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__1_ccff_tail),
    .chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__25_ccff_tail)
  );


  cbx_1__1_
  cbx_3__11_
  (
    .clk_1_S_out(clk_1_wires[81]),
    .clk_1_N_out(clk_1_wires[80]),
    .clk_1_E_in(clk_1_wires[79]),
    .prog_clk_1_S_out(prog_clk_1_wires[81]),
    .prog_clk_1_N_out(prog_clk_1_wires[80]),
    .prog_clk_1_E_in(prog_clk_1_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[134]),
    .config_enable_S_out(config_enableWires[562]),
    .config_enable_E_in(config_enableWires[561]),
    .config_enable_W_out(config_enableWires[560]),
    .sc_head_S_out(sc_headWires[56]),
    .sc_head_N_in(sc_headWires[55]),
    .pReset_S_out(pResetWires[562]),
    .pReset_E_in(pResetWires[561]),
    .pReset_W_out(pResetWires[560]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[32]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[32]),
    .chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__13_ccff_tail),
    .chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__26_ccff_tail)
  );


  cbx_1__1_
  cbx_4__1_
  (
    .clk_1_S_out(clk_1_wires[48]),
    .clk_1_N_out(clk_1_wires[47]),
    .clk_1_W_in(clk_1_wires[43]),
    .prog_clk_1_S_out(prog_clk_1_wires[48]),
    .prog_clk_1_N_out(prog_clk_1_wires[47]),
    .prog_clk_1_W_in(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[142]),
    .config_enable_S_out(config_enableWires[76]),
    .config_enable_E_in(config_enableWires[75]),
    .config_enable_W_out(config_enableWires[74]),
    .sc_head_N_out(sc_headWires[82]),
    .sc_head_S_in(sc_headWires[81]),
    .pReset_S_out(pResetWires[76]),
    .pReset_E_in(pResetWires[75]),
    .pReset_W_out(pResetWires[74]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[33]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[33]),
    .chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__14_ccff_tail),
    .chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__27_ccff_tail)
  );


  cbx_1__1_
  cbx_4__2_
  (
    .clk_2_W_out(clk_2_wires[28]),
    .clk_2_E_in(clk_2_wires[27]),
    .prog_clk_2_W_out(prog_clk_2_wires[28]),
    .prog_clk_2_E_in(prog_clk_2_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[145]),
    .config_enable_S_out(config_enableWires[125]),
    .config_enable_E_in(config_enableWires[124]),
    .config_enable_W_out(config_enableWires[123]),
    .sc_head_N_out(sc_headWires[84]),
    .sc_head_S_in(sc_headWires[83]),
    .pReset_S_out(pResetWires[125]),
    .pReset_E_in(pResetWires[124]),
    .pReset_W_out(pResetWires[123]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[34]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[34]),
    .chanx_left_in(sb_1__2__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__2_ccff_tail),
    .chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__28_ccff_tail)
  );


  cbx_1__1_
  cbx_4__4_
  (
    .clk_2_W_out(clk_2_wires[37]),
    .clk_2_E_in(clk_2_wires[36]),
    .prog_clk_2_W_out(prog_clk_2_wires[37]),
    .prog_clk_2_E_in(prog_clk_2_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[151]),
    .config_enable_S_out(config_enableWires[223]),
    .config_enable_E_in(config_enableWires[222]),
    .config_enable_W_out(config_enableWires[221]),
    .sc_head_N_out(sc_headWires[88]),
    .sc_head_S_in(sc_headWires[87]),
    .pReset_S_out(pResetWires[223]),
    .pReset_E_in(pResetWires[222]),
    .pReset_W_out(pResetWires[221]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[36]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[36]),
    .chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__15_ccff_tail),
    .chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__29_ccff_tail)
  );


  cbx_1__1_
  cbx_4__5_
  (
    .clk_1_S_out(clk_1_wires[62]),
    .clk_1_N_out(clk_1_wires[61]),
    .clk_1_W_in(clk_1_wires[57]),
    .prog_clk_1_S_out(prog_clk_1_wires[62]),
    .prog_clk_1_N_out(prog_clk_1_wires[61]),
    .prog_clk_1_W_in(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[154]),
    .config_enable_S_out(config_enableWires[272]),
    .config_enable_E_in(config_enableWires[271]),
    .config_enable_W_out(config_enableWires[270]),
    .sc_head_N_out(sc_headWires[90]),
    .sc_head_S_in(sc_headWires[89]),
    .pReset_S_out(pResetWires[272]),
    .pReset_E_in(pResetWires[271]),
    .pReset_W_out(pResetWires[270]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[37]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[37]),
    .chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__16_ccff_tail),
    .chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__30_ccff_tail)
  );


  cbx_1__1_
  cbx_4__6_
  (
    .clk_3_W_out(clk_3_wires[47]),
    .clk_3_E_in(clk_3_wires[46]),
    .prog_clk_3_W_out(prog_clk_3_wires[47]),
    .prog_clk_3_E_in(prog_clk_3_wires[46]),
    .prog_clk_0_N_in(prog_clk_0_wires[157]),
    .config_enable_S_out(config_enableWires[321]),
    .config_enable_E_in(config_enableWires[320]),
    .config_enable_W_out(config_enableWires[319]),
    .sc_head_N_out(sc_headWires[92]),
    .sc_head_S_in(sc_headWires[91]),
    .pReset_S_out(pResetWires[321]),
    .pReset_E_in(pResetWires[320]),
    .pReset_W_out(pResetWires[319]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[38]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[38]),
    .chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__17_ccff_tail),
    .chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__31_ccff_tail)
  );


  cbx_1__1_
  cbx_4__7_
  (
    .clk_1_S_out(clk_1_wires[69]),
    .clk_1_N_out(clk_1_wires[68]),
    .clk_1_W_in(clk_1_wires[64]),
    .prog_clk_1_S_out(prog_clk_1_wires[69]),
    .prog_clk_1_N_out(prog_clk_1_wires[68]),
    .prog_clk_1_W_in(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[160]),
    .config_enable_S_out(config_enableWires[370]),
    .config_enable_E_in(config_enableWires[369]),
    .config_enable_W_out(config_enableWires[368]),
    .sc_head_N_out(sc_headWires[94]),
    .sc_head_S_in(sc_headWires[93]),
    .pReset_S_out(pResetWires[370]),
    .pReset_E_in(pResetWires[369]),
    .pReset_W_out(pResetWires[368]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[39]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[39]),
    .chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__18_ccff_tail),
    .chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__32_ccff_tail)
  );


  cbx_1__1_
  cbx_4__8_
  (
    .clk_2_W_out(clk_2_wires[50]),
    .clk_2_E_in(clk_2_wires[49]),
    .prog_clk_2_W_out(prog_clk_2_wires[50]),
    .prog_clk_2_E_in(prog_clk_2_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[163]),
    .config_enable_S_out(config_enableWires[419]),
    .config_enable_E_in(config_enableWires[418]),
    .config_enable_W_out(config_enableWires[417]),
    .sc_head_N_out(sc_headWires[96]),
    .sc_head_S_in(sc_headWires[95]),
    .pReset_S_out(pResetWires[419]),
    .pReset_E_in(pResetWires[418]),
    .pReset_W_out(pResetWires[417]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[40]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[40]),
    .chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__19_ccff_tail),
    .chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__33_ccff_tail)
  );


  cbx_1__1_
  cbx_4__9_
  (
    .clk_1_S_out(clk_1_wires[76]),
    .clk_1_N_out(clk_1_wires[75]),
    .clk_1_W_in(clk_1_wires[71]),
    .prog_clk_1_S_out(prog_clk_1_wires[76]),
    .prog_clk_1_N_out(prog_clk_1_wires[75]),
    .prog_clk_1_W_in(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[166]),
    .config_enable_S_out(config_enableWires[468]),
    .config_enable_E_in(config_enableWires[467]),
    .config_enable_W_out(config_enableWires[466]),
    .sc_head_N_out(sc_headWires[98]),
    .sc_head_S_in(sc_headWires[97]),
    .pReset_S_out(pResetWires[468]),
    .pReset_E_in(pResetWires[467]),
    .pReset_W_out(pResetWires[466]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[41]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[41]),
    .chanx_left_in(sb_1__2__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__3_ccff_tail),
    .chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__34_ccff_tail)
  );


  cbx_1__1_
  cbx_4__11_
  (
    .clk_1_S_out(clk_1_wires[83]),
    .clk_1_N_out(clk_1_wires[82]),
    .clk_1_W_in(clk_1_wires[78]),
    .prog_clk_1_S_out(prog_clk_1_wires[83]),
    .prog_clk_1_N_out(prog_clk_1_wires[82]),
    .prog_clk_1_W_in(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[172]),
    .config_enable_S_out(config_enableWires[566]),
    .config_enable_E_in(config_enableWires[565]),
    .config_enable_W_out(config_enableWires[564]),
    .sc_head_N_out(sc_headWires[102]),
    .sc_head_S_in(sc_headWires[101]),
    .pReset_S_out(pResetWires[566]),
    .pReset_E_in(pResetWires[565]),
    .pReset_W_out(pResetWires[564]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[43]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[43]),
    .chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__20_ccff_tail),
    .chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__35_ccff_tail)
  );


  cbx_1__1_
  cbx_5__1_
  (
    .clk_1_S_out(clk_1_wires[88]),
    .clk_1_N_out(clk_1_wires[87]),
    .clk_1_E_in(clk_1_wires[86]),
    .prog_clk_1_S_out(prog_clk_1_wires[88]),
    .prog_clk_1_N_out(prog_clk_1_wires[87]),
    .prog_clk_1_E_in(prog_clk_1_wires[86]),
    .prog_clk_0_N_in(prog_clk_0_wires[180]),
    .config_enable_S_out(config_enableWires[80]),
    .config_enable_E_in(config_enableWires[79]),
    .config_enable_W_out(config_enableWires[78]),
    .sc_head_S_out(sc_headWires[128]),
    .sc_head_N_in(sc_headWires[127]),
    .pReset_S_out(pResetWires[80]),
    .pReset_E_in(pResetWires[79]),
    .pReset_W_out(pResetWires[78]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[44]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[44]),
    .chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__21_ccff_tail),
    .chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__36_ccff_tail)
  );


  cbx_1__1_
  cbx_5__2_
  (
    .clk_2_E_out(clk_2_wires[26]),
    .clk_2_W_in(clk_2_wires[25]),
    .prog_clk_2_E_out(prog_clk_2_wires[26]),
    .prog_clk_2_W_in(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[183]),
    .config_enable_S_out(config_enableWires[129]),
    .config_enable_E_in(config_enableWires[128]),
    .config_enable_W_out(config_enableWires[127]),
    .sc_head_S_out(sc_headWires[126]),
    .sc_head_N_in(sc_headWires[125]),
    .pReset_S_out(pResetWires[129]),
    .pReset_E_in(pResetWires[128]),
    .pReset_W_out(pResetWires[127]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[45]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[45]),
    .chanx_left_in(sb_2__2__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__4_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__2_ccff_tail),
    .chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__37_ccff_tail)
  );


  cbx_1__1_
  cbx_5__4_
  (
    .clk_2_E_out(clk_2_wires[35]),
    .clk_2_W_in(clk_2_wires[34]),
    .prog_clk_2_E_out(prog_clk_2_wires[35]),
    .prog_clk_2_W_in(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[189]),
    .config_enable_S_out(config_enableWires[227]),
    .config_enable_E_in(config_enableWires[226]),
    .config_enable_W_out(config_enableWires[225]),
    .sc_head_S_out(sc_headWires[122]),
    .sc_head_N_in(sc_headWires[121]),
    .pReset_S_out(pResetWires[227]),
    .pReset_E_in(pResetWires[226]),
    .pReset_W_out(pResetWires[225]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[47]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[47]),
    .chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__22_ccff_tail),
    .chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__38_ccff_tail)
  );


  cbx_1__1_
  cbx_5__5_
  (
    .clk_1_S_out(clk_1_wires[102]),
    .clk_1_N_out(clk_1_wires[101]),
    .clk_1_E_in(clk_1_wires[100]),
    .prog_clk_1_S_out(prog_clk_1_wires[102]),
    .prog_clk_1_N_out(prog_clk_1_wires[101]),
    .prog_clk_1_E_in(prog_clk_1_wires[100]),
    .prog_clk_0_N_in(prog_clk_0_wires[192]),
    .config_enable_S_out(config_enableWires[276]),
    .config_enable_E_in(config_enableWires[275]),
    .config_enable_W_out(config_enableWires[274]),
    .sc_head_S_out(sc_headWires[120]),
    .sc_head_N_in(sc_headWires[119]),
    .pReset_S_out(pResetWires[276]),
    .pReset_E_in(pResetWires[275]),
    .pReset_W_out(pResetWires[274]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[48]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[48]),
    .chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__23_ccff_tail),
    .chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__39_ccff_tail)
  );


  cbx_1__1_
  cbx_5__6_
  (
    .clk_3_W_out(clk_3_wires[7]),
    .clk_3_E_in(clk_3_wires[6]),
    .prog_clk_3_W_out(prog_clk_3_wires[7]),
    .prog_clk_3_E_in(prog_clk_3_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[195]),
    .config_enable_S_out(config_enableWires[325]),
    .config_enable_E_in(config_enableWires[324]),
    .config_enable_W_out(config_enableWires[323]),
    .sc_head_S_out(sc_headWires[118]),
    .sc_head_N_in(sc_headWires[117]),
    .pReset_S_out(pResetWires[325]),
    .pReset_E_in(pResetWires[324]),
    .pReset_W_out(pResetWires[323]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[49]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[49]),
    .chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__24_ccff_tail),
    .chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__40_ccff_tail)
  );


  cbx_1__1_
  cbx_5__7_
  (
    .clk_1_S_out(clk_1_wires[109]),
    .clk_1_N_out(clk_1_wires[108]),
    .clk_1_E_in(clk_1_wires[107]),
    .prog_clk_1_S_out(prog_clk_1_wires[109]),
    .prog_clk_1_N_out(prog_clk_1_wires[108]),
    .prog_clk_1_E_in(prog_clk_1_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[198]),
    .config_enable_S_out(config_enableWires[374]),
    .config_enable_E_in(config_enableWires[373]),
    .config_enable_W_out(config_enableWires[372]),
    .sc_head_S_out(sc_headWires[116]),
    .sc_head_N_in(sc_headWires[115]),
    .pReset_S_out(pResetWires[374]),
    .pReset_E_in(pResetWires[373]),
    .pReset_W_out(pResetWires[372]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[50]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[50]),
    .chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__25_ccff_tail),
    .chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__41_ccff_tail)
  );


  cbx_1__1_
  cbx_5__8_
  (
    .clk_2_E_out(clk_2_wires[48]),
    .clk_2_W_in(clk_2_wires[47]),
    .prog_clk_2_E_out(prog_clk_2_wires[48]),
    .prog_clk_2_W_in(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[201]),
    .config_enable_S_out(config_enableWires[423]),
    .config_enable_E_in(config_enableWires[422]),
    .config_enable_W_out(config_enableWires[421]),
    .sc_head_S_out(sc_headWires[114]),
    .sc_head_N_in(sc_headWires[113]),
    .pReset_S_out(pResetWires[423]),
    .pReset_E_in(pResetWires[422]),
    .pReset_W_out(pResetWires[421]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[51]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[51]),
    .chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__26_ccff_tail),
    .chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__42_ccff_tail)
  );


  cbx_1__1_
  cbx_5__9_
  (
    .clk_1_S_out(clk_1_wires[116]),
    .clk_1_N_out(clk_1_wires[115]),
    .clk_1_E_in(clk_1_wires[114]),
    .prog_clk_1_S_out(prog_clk_1_wires[116]),
    .prog_clk_1_N_out(prog_clk_1_wires[115]),
    .prog_clk_1_E_in(prog_clk_1_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[204]),
    .config_enable_S_out(config_enableWires[472]),
    .config_enable_E_in(config_enableWires[471]),
    .config_enable_W_out(config_enableWires[470]),
    .sc_head_S_out(sc_headWires[112]),
    .sc_head_N_in(sc_headWires[111]),
    .pReset_S_out(pResetWires[472]),
    .pReset_E_in(pResetWires[471]),
    .pReset_W_out(pResetWires[470]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[52]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[52]),
    .chanx_left_in(sb_2__2__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__5_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__3_ccff_tail),
    .chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__43_ccff_tail)
  );


  cbx_1__1_
  cbx_5__11_
  (
    .clk_1_S_out(clk_1_wires[123]),
    .clk_1_N_out(clk_1_wires[122]),
    .clk_1_E_in(clk_1_wires[121]),
    .prog_clk_1_S_out(prog_clk_1_wires[123]),
    .prog_clk_1_N_out(prog_clk_1_wires[122]),
    .prog_clk_1_E_in(prog_clk_1_wires[121]),
    .prog_clk_0_N_in(prog_clk_0_wires[210]),
    .config_enable_S_out(config_enableWires[570]),
    .config_enable_E_in(config_enableWires[569]),
    .config_enable_W_out(config_enableWires[568]),
    .sc_head_S_out(sc_headWires[108]),
    .sc_head_N_in(sc_headWires[107]),
    .pReset_S_out(pResetWires[570]),
    .pReset_E_in(pResetWires[569]),
    .pReset_W_out(pResetWires[568]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[54]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[54]),
    .chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__27_ccff_tail),
    .chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__44_ccff_tail)
  );


  cbx_1__1_
  cbx_6__1_
  (
    .clk_1_S_out(clk_1_wires[90]),
    .clk_1_N_out(clk_1_wires[89]),
    .clk_1_W_in(clk_1_wires[85]),
    .prog_clk_1_S_out(prog_clk_1_wires[90]),
    .prog_clk_1_N_out(prog_clk_1_wires[89]),
    .prog_clk_1_W_in(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[218]),
    .config_enable_S_out(config_enableWires[84]),
    .config_enable_E_in(config_enableWires[83]),
    .config_enable_W_out(config_enableWires[82]),
    .sc_head_N_out(sc_headWires[134]),
    .sc_head_S_in(sc_headWires[133]),
    .pReset_S_out(pResetWires[84]),
    .pReset_E_in(pResetWires[83]),
    .pReset_W_out(pResetWires[82]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[55]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[55]),
    .chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__28_ccff_tail),
    .chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__45_ccff_tail)
  );


  cbx_1__1_
  cbx_6__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[221]),
    .config_enable_S_out(config_enableWires[133]),
    .config_enable_E_in(config_enableWires[132]),
    .config_enable_W_out(config_enableWires[131]),
    .sc_head_N_out(sc_headWires[136]),
    .sc_head_S_in(sc_headWires[135]),
    .pReset_S_out(pResetWires[133]),
    .pReset_E_in(pResetWires[132]),
    .pReset_W_out(pResetWires[131]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[56]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[56]),
    .chanx_left_in(sb_1__2__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__4_ccff_tail),
    .chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__46_ccff_tail)
  );


  cbx_1__1_
  cbx_6__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[227]),
    .config_enable_S_out(config_enableWires[231]),
    .config_enable_E_in(config_enableWires[230]),
    .config_enable_W_out(config_enableWires[229]),
    .sc_head_N_out(sc_headWires[140]),
    .sc_head_S_in(sc_headWires[139]),
    .pReset_S_out(pResetWires[231]),
    .pReset_E_in(pResetWires[230]),
    .pReset_W_out(pResetWires[229]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[58]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[58]),
    .chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__29_ccff_tail),
    .chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__47_ccff_tail)
  );


  cbx_1__1_
  cbx_6__5_
  (
    .clk_1_S_out(clk_1_wires[104]),
    .clk_1_N_out(clk_1_wires[103]),
    .clk_1_W_in(clk_1_wires[99]),
    .prog_clk_1_S_out(prog_clk_1_wires[104]),
    .prog_clk_1_N_out(prog_clk_1_wires[103]),
    .prog_clk_1_W_in(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[230]),
    .config_enable_S_out(config_enableWires[280]),
    .config_enable_E_in(config_enableWires[279]),
    .config_enable_W_out(config_enableWires[278]),
    .sc_head_N_out(sc_headWires[142]),
    .sc_head_S_in(sc_headWires[141]),
    .pReset_S_out(pResetWires[280]),
    .pReset_E_in(pResetWires[279]),
    .pReset_W_out(pResetWires[278]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[59]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[59]),
    .chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__30_ccff_tail),
    .chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__48_ccff_tail)
  );


  cbx_1__1_
  cbx_6__6_
  (
    .clk_3_W_out(clk_3_wires[3]),
    .clk_3_E_in(clk_3_wires[2]),
    .prog_clk_3_W_out(prog_clk_3_wires[3]),
    .prog_clk_3_E_in(prog_clk_3_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[233]),
    .config_enable_S_out(config_enableWires[329]),
    .config_enable_E_in(config_enableWires[328]),
    .config_enable_W_out(config_enableWires[327]),
    .sc_head_N_out(sc_headWires[144]),
    .sc_head_S_in(sc_headWires[143]),
    .pReset_S_out(pResetWires[329]),
    .pReset_E_in(pResetWires[328]),
    .pReset_W_out(pResetWires[327]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[60]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[60]),
    .chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__31_ccff_tail),
    .chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__49_ccff_tail)
  );


  cbx_1__1_
  cbx_6__7_
  (
    .clk_1_S_out(clk_1_wires[111]),
    .clk_1_N_out(clk_1_wires[110]),
    .clk_1_W_in(clk_1_wires[106]),
    .prog_clk_1_S_out(prog_clk_1_wires[111]),
    .prog_clk_1_N_out(prog_clk_1_wires[110]),
    .prog_clk_1_W_in(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[236]),
    .config_enable_S_out(config_enableWires[378]),
    .config_enable_E_in(config_enableWires[377]),
    .config_enable_W_out(config_enableWires[376]),
    .sc_head_N_out(sc_headWires[146]),
    .sc_head_S_in(sc_headWires[145]),
    .pReset_S_out(pResetWires[378]),
    .pReset_E_in(pResetWires[377]),
    .pReset_W_out(pResetWires[376]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[61]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[61]),
    .chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__32_ccff_tail),
    .chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__50_ccff_tail)
  );


  cbx_1__1_
  cbx_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[239]),
    .config_enable_S_out(config_enableWires[427]),
    .config_enable_E_in(config_enableWires[426]),
    .config_enable_W_out(config_enableWires[425]),
    .sc_head_N_out(sc_headWires[148]),
    .sc_head_S_in(sc_headWires[147]),
    .pReset_S_out(pResetWires[427]),
    .pReset_E_in(pResetWires[426]),
    .pReset_W_out(pResetWires[425]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[62]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[62]),
    .chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__33_ccff_tail),
    .chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__51_ccff_tail)
  );


  cbx_1__1_
  cbx_6__9_
  (
    .clk_1_S_out(clk_1_wires[118]),
    .clk_1_N_out(clk_1_wires[117]),
    .clk_1_W_in(clk_1_wires[113]),
    .prog_clk_1_S_out(prog_clk_1_wires[118]),
    .prog_clk_1_N_out(prog_clk_1_wires[117]),
    .prog_clk_1_W_in(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[242]),
    .config_enable_S_out(config_enableWires[476]),
    .config_enable_E_in(config_enableWires[475]),
    .config_enable_W_out(config_enableWires[474]),
    .sc_head_N_out(sc_headWires[150]),
    .sc_head_S_in(sc_headWires[149]),
    .pReset_S_out(pResetWires[476]),
    .pReset_E_in(pResetWires[475]),
    .pReset_W_out(pResetWires[474]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[63]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[63]),
    .chanx_left_in(sb_1__2__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__5_ccff_tail),
    .chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__52_ccff_tail)
  );


  cbx_1__1_
  cbx_6__11_
  (
    .clk_1_S_out(clk_1_wires[125]),
    .clk_1_N_out(clk_1_wires[124]),
    .clk_1_W_in(clk_1_wires[120]),
    .prog_clk_1_S_out(prog_clk_1_wires[125]),
    .prog_clk_1_N_out(prog_clk_1_wires[124]),
    .prog_clk_1_W_in(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[248]),
    .config_enable_S_out(config_enableWires[574]),
    .config_enable_E_in(config_enableWires[573]),
    .config_enable_W_out(config_enableWires[572]),
    .sc_head_N_out(sc_headWires[154]),
    .sc_head_S_in(sc_headWires[153]),
    .pReset_S_out(pResetWires[574]),
    .pReset_E_in(pResetWires[573]),
    .pReset_W_out(pResetWires[572]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[65]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[65]),
    .chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__34_ccff_tail),
    .chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__53_ccff_tail)
  );


  cbx_1__1_
  cbx_7__1_
  (
    .clk_1_S_out(clk_1_wires[130]),
    .clk_1_N_out(clk_1_wires[129]),
    .clk_1_E_in(clk_1_wires[128]),
    .prog_clk_1_S_out(prog_clk_1_wires[130]),
    .prog_clk_1_N_out(prog_clk_1_wires[129]),
    .prog_clk_1_E_in(prog_clk_1_wires[128]),
    .prog_clk_0_N_in(prog_clk_0_wires[256]),
    .config_enable_S_out(config_enableWires[88]),
    .config_enable_E_out(config_enableWires[87]),
    .config_enable_W_in(config_enableWires[86]),
    .sc_head_S_out(sc_headWires[180]),
    .sc_head_N_in(sc_headWires[179]),
    .pReset_S_out(pResetWires[88]),
    .pReset_E_out(pResetWires[87]),
    .pReset_W_in(pResetWires[86]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[66]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[66]),
    .chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__35_ccff_tail),
    .chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__54_ccff_tail)
  );


  cbx_1__1_
  cbx_7__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[259]),
    .config_enable_S_out(config_enableWires[137]),
    .config_enable_E_out(config_enableWires[136]),
    .config_enable_W_in(config_enableWires[135]),
    .sc_head_S_out(sc_headWires[178]),
    .sc_head_N_in(sc_headWires[177]),
    .pReset_S_out(pResetWires[137]),
    .pReset_E_out(pResetWires[136]),
    .pReset_W_in(pResetWires[135]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[67]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[67]),
    .chanx_left_in(sb_2__2__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__6_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__4_ccff_tail),
    .chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__55_ccff_tail)
  );


  cbx_1__1_
  cbx_7__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[265]),
    .config_enable_S_out(config_enableWires[235]),
    .config_enable_E_out(config_enableWires[234]),
    .config_enable_W_in(config_enableWires[233]),
    .sc_head_S_out(sc_headWires[174]),
    .sc_head_N_in(sc_headWires[173]),
    .pReset_S_out(pResetWires[235]),
    .pReset_E_out(pResetWires[234]),
    .pReset_W_in(pResetWires[233]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[69]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[69]),
    .chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__36_ccff_tail),
    .chanx_left_out(cbx_1__1__56_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__56_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__56_ccff_tail)
  );


  cbx_1__1_
  cbx_7__5_
  (
    .clk_1_S_out(clk_1_wires[144]),
    .clk_1_N_out(clk_1_wires[143]),
    .clk_1_E_in(clk_1_wires[142]),
    .prog_clk_1_S_out(prog_clk_1_wires[144]),
    .prog_clk_1_N_out(prog_clk_1_wires[143]),
    .prog_clk_1_E_in(prog_clk_1_wires[142]),
    .prog_clk_0_N_in(prog_clk_0_wires[268]),
    .config_enable_S_out(config_enableWires[284]),
    .config_enable_E_out(config_enableWires[283]),
    .config_enable_W_in(config_enableWires[282]),
    .sc_head_S_out(sc_headWires[172]),
    .sc_head_N_in(sc_headWires[171]),
    .pReset_S_out(pResetWires[284]),
    .pReset_E_out(pResetWires[283]),
    .pReset_W_in(pResetWires[282]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[70]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[70]),
    .chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__37_ccff_tail),
    .chanx_left_out(cbx_1__1__57_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__57_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__57_ccff_tail)
  );


  cbx_1__1_
  cbx_7__6_
  (
    .clk_3_E_out(clk_3_wires[1]),
    .clk_3_W_in(clk_3_wires[0]),
    .prog_clk_3_E_out(prog_clk_3_wires[1]),
    .prog_clk_3_W_in(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[271]),
    .config_enable_S_out(config_enableWires[333]),
    .config_enable_E_out(config_enableWires[332]),
    .config_enable_W_in(config_enableWires[331]),
    .sc_head_S_out(sc_headWires[170]),
    .sc_head_N_in(sc_headWires[169]),
    .pReset_S_out(pResetWires[333]),
    .pReset_E_out(pResetWires[332]),
    .pReset_W_in(pResetWires[331]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[71]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[71]),
    .chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__38_ccff_tail),
    .chanx_left_out(cbx_1__1__58_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__58_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__58_ccff_tail)
  );


  cbx_1__1_
  cbx_7__7_
  (
    .clk_1_S_out(clk_1_wires[151]),
    .clk_1_N_out(clk_1_wires[150]),
    .clk_1_E_in(clk_1_wires[149]),
    .prog_clk_1_S_out(prog_clk_1_wires[151]),
    .prog_clk_1_N_out(prog_clk_1_wires[150]),
    .prog_clk_1_E_in(prog_clk_1_wires[149]),
    .prog_clk_0_N_in(prog_clk_0_wires[274]),
    .config_enable_S_out(config_enableWires[382]),
    .config_enable_E_out(config_enableWires[381]),
    .config_enable_W_in(config_enableWires[380]),
    .sc_head_S_out(sc_headWires[168]),
    .sc_head_N_in(sc_headWires[167]),
    .pReset_S_out(pResetWires[382]),
    .pReset_E_out(pResetWires[381]),
    .pReset_W_in(pResetWires[380]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[72]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[72]),
    .chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__39_ccff_tail),
    .chanx_left_out(cbx_1__1__59_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__59_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__59_ccff_tail)
  );


  cbx_1__1_
  cbx_7__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[277]),
    .config_enable_S_out(config_enableWires[431]),
    .config_enable_E_out(config_enableWires[430]),
    .config_enable_W_in(config_enableWires[429]),
    .sc_head_S_out(sc_headWires[166]),
    .sc_head_N_in(sc_headWires[165]),
    .pReset_S_out(pResetWires[431]),
    .pReset_E_out(pResetWires[430]),
    .pReset_W_in(pResetWires[429]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[73]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[73]),
    .chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__40_ccff_tail),
    .chanx_left_out(cbx_1__1__60_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__60_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__60_ccff_tail)
  );


  cbx_1__1_
  cbx_7__9_
  (
    .clk_1_S_out(clk_1_wires[158]),
    .clk_1_N_out(clk_1_wires[157]),
    .clk_1_E_in(clk_1_wires[156]),
    .prog_clk_1_S_out(prog_clk_1_wires[158]),
    .prog_clk_1_N_out(prog_clk_1_wires[157]),
    .prog_clk_1_E_in(prog_clk_1_wires[156]),
    .prog_clk_0_N_in(prog_clk_0_wires[280]),
    .config_enable_S_out(config_enableWires[480]),
    .config_enable_E_out(config_enableWires[479]),
    .config_enable_W_in(config_enableWires[478]),
    .sc_head_S_out(sc_headWires[164]),
    .sc_head_N_in(sc_headWires[163]),
    .pReset_S_out(pResetWires[480]),
    .pReset_E_out(pResetWires[479]),
    .pReset_W_in(pResetWires[478]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[74]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[74]),
    .chanx_left_in(sb_2__2__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__7_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__5_ccff_tail),
    .chanx_left_out(cbx_1__1__61_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__61_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__61_ccff_tail)
  );


  cbx_1__1_
  cbx_7__11_
  (
    .clk_1_S_out(clk_1_wires[165]),
    .clk_1_N_out(clk_1_wires[164]),
    .clk_1_E_in(clk_1_wires[163]),
    .prog_clk_1_S_out(prog_clk_1_wires[165]),
    .prog_clk_1_N_out(prog_clk_1_wires[164]),
    .prog_clk_1_E_in(prog_clk_1_wires[163]),
    .prog_clk_0_N_in(prog_clk_0_wires[286]),
    .config_enable_S_out(config_enableWires[578]),
    .config_enable_E_out(config_enableWires[577]),
    .config_enable_W_in(config_enableWires[576]),
    .sc_head_S_out(sc_headWires[160]),
    .sc_head_N_in(sc_headWires[159]),
    .pReset_S_out(pResetWires[578]),
    .pReset_E_out(pResetWires[577]),
    .pReset_W_in(pResetWires[576]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[76]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[76]),
    .chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__41_ccff_tail),
    .chanx_left_out(cbx_1__1__62_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__62_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__62_ccff_tail)
  );


  cbx_1__1_
  cbx_8__1_
  (
    .clk_1_S_out(clk_1_wires[132]),
    .clk_1_N_out(clk_1_wires[131]),
    .clk_1_W_in(clk_1_wires[127]),
    .prog_clk_1_S_out(prog_clk_1_wires[132]),
    .prog_clk_1_N_out(prog_clk_1_wires[131]),
    .prog_clk_1_W_in(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[294]),
    .config_enable_S_out(config_enableWires[92]),
    .config_enable_E_out(config_enableWires[91]),
    .config_enable_W_in(config_enableWires[90]),
    .sc_head_N_out(sc_headWires[186]),
    .sc_head_S_in(sc_headWires[185]),
    .pReset_S_out(pResetWires[92]),
    .pReset_E_out(pResetWires[91]),
    .pReset_W_in(pResetWires[90]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[77]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[77]),
    .chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__42_ccff_tail),
    .chanx_left_out(cbx_1__1__63_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__63_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__63_ccff_tail)
  );


  cbx_1__1_
  cbx_8__2_
  (
    .clk_2_W_out(clk_2_wires[72]),
    .clk_2_E_in(clk_2_wires[71]),
    .prog_clk_2_W_out(prog_clk_2_wires[72]),
    .prog_clk_2_E_in(prog_clk_2_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[297]),
    .config_enable_S_out(config_enableWires[141]),
    .config_enable_E_out(config_enableWires[140]),
    .config_enable_W_in(config_enableWires[139]),
    .sc_head_N_out(sc_headWires[188]),
    .sc_head_S_in(sc_headWires[187]),
    .pReset_S_out(pResetWires[141]),
    .pReset_E_out(pResetWires[140]),
    .pReset_W_in(pResetWires[139]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[78]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[78]),
    .chanx_left_in(sb_1__2__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__6_ccff_tail),
    .chanx_left_out(cbx_1__1__64_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__64_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__64_ccff_tail)
  );


  cbx_1__1_
  cbx_8__4_
  (
    .clk_2_W_out(clk_2_wires[81]),
    .clk_2_E_in(clk_2_wires[80]),
    .prog_clk_2_W_out(prog_clk_2_wires[81]),
    .prog_clk_2_E_in(prog_clk_2_wires[80]),
    .prog_clk_0_N_in(prog_clk_0_wires[303]),
    .config_enable_S_out(config_enableWires[239]),
    .config_enable_E_out(config_enableWires[238]),
    .config_enable_W_in(config_enableWires[237]),
    .sc_head_N_out(sc_headWires[192]),
    .sc_head_S_in(sc_headWires[191]),
    .pReset_S_out(pResetWires[239]),
    .pReset_E_out(pResetWires[238]),
    .pReset_W_in(pResetWires[237]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[80]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[80]),
    .chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__43_ccff_tail),
    .chanx_left_out(cbx_1__1__65_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__65_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__65_ccff_tail)
  );


  cbx_1__1_
  cbx_8__5_
  (
    .clk_1_S_out(clk_1_wires[146]),
    .clk_1_N_out(clk_1_wires[145]),
    .clk_1_W_in(clk_1_wires[141]),
    .prog_clk_1_S_out(prog_clk_1_wires[146]),
    .prog_clk_1_N_out(prog_clk_1_wires[145]),
    .prog_clk_1_W_in(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[306]),
    .config_enable_S_out(config_enableWires[288]),
    .config_enable_E_out(config_enableWires[287]),
    .config_enable_W_in(config_enableWires[286]),
    .sc_head_N_out(sc_headWires[194]),
    .sc_head_S_in(sc_headWires[193]),
    .pReset_S_out(pResetWires[288]),
    .pReset_E_out(pResetWires[287]),
    .pReset_W_in(pResetWires[286]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[81]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[81]),
    .chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__44_ccff_tail),
    .chanx_left_out(cbx_1__1__66_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__66_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__66_ccff_tail)
  );


  cbx_1__1_
  cbx_8__6_
  (
    .clk_3_E_out(clk_3_wires[5]),
    .clk_3_W_in(clk_3_wires[4]),
    .prog_clk_3_E_out(prog_clk_3_wires[5]),
    .prog_clk_3_W_in(prog_clk_3_wires[4]),
    .prog_clk_0_N_in(prog_clk_0_wires[309]),
    .config_enable_S_out(config_enableWires[337]),
    .config_enable_E_out(config_enableWires[336]),
    .config_enable_W_in(config_enableWires[335]),
    .sc_head_N_out(sc_headWires[196]),
    .sc_head_S_in(sc_headWires[195]),
    .pReset_S_out(pResetWires[337]),
    .pReset_E_out(pResetWires[336]),
    .pReset_W_in(pResetWires[335]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[82]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[82]),
    .chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__45_ccff_tail),
    .chanx_left_out(cbx_1__1__67_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__67_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__67_ccff_tail)
  );


  cbx_1__1_
  cbx_8__7_
  (
    .clk_1_S_out(clk_1_wires[153]),
    .clk_1_N_out(clk_1_wires[152]),
    .clk_1_W_in(clk_1_wires[148]),
    .prog_clk_1_S_out(prog_clk_1_wires[153]),
    .prog_clk_1_N_out(prog_clk_1_wires[152]),
    .prog_clk_1_W_in(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[312]),
    .config_enable_S_out(config_enableWires[386]),
    .config_enable_E_out(config_enableWires[385]),
    .config_enable_W_in(config_enableWires[384]),
    .sc_head_N_out(sc_headWires[198]),
    .sc_head_S_in(sc_headWires[197]),
    .pReset_S_out(pResetWires[386]),
    .pReset_E_out(pResetWires[385]),
    .pReset_W_in(pResetWires[384]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[83]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[83]),
    .chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__46_ccff_tail),
    .chanx_left_out(cbx_1__1__68_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__68_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__68_ccff_tail)
  );


  cbx_1__1_
  cbx_8__8_
  (
    .clk_2_W_out(clk_2_wires[94]),
    .clk_2_E_in(clk_2_wires[93]),
    .prog_clk_2_W_out(prog_clk_2_wires[94]),
    .prog_clk_2_E_in(prog_clk_2_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[315]),
    .config_enable_S_out(config_enableWires[435]),
    .config_enable_E_out(config_enableWires[434]),
    .config_enable_W_in(config_enableWires[433]),
    .sc_head_N_out(sc_headWires[200]),
    .sc_head_S_in(sc_headWires[199]),
    .pReset_S_out(pResetWires[435]),
    .pReset_E_out(pResetWires[434]),
    .pReset_W_in(pResetWires[433]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[84]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[84]),
    .chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__47_ccff_tail),
    .chanx_left_out(cbx_1__1__69_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__69_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__69_ccff_tail)
  );


  cbx_1__1_
  cbx_8__9_
  (
    .clk_1_S_out(clk_1_wires[160]),
    .clk_1_N_out(clk_1_wires[159]),
    .clk_1_W_in(clk_1_wires[155]),
    .prog_clk_1_S_out(prog_clk_1_wires[160]),
    .prog_clk_1_N_out(prog_clk_1_wires[159]),
    .prog_clk_1_W_in(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[318]),
    .config_enable_S_out(config_enableWires[484]),
    .config_enable_E_out(config_enableWires[483]),
    .config_enable_W_in(config_enableWires[482]),
    .sc_head_N_out(sc_headWires[202]),
    .sc_head_S_in(sc_headWires[201]),
    .pReset_S_out(pResetWires[484]),
    .pReset_E_out(pResetWires[483]),
    .pReset_W_in(pResetWires[482]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[85]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[85]),
    .chanx_left_in(sb_1__2__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__7_ccff_tail),
    .chanx_left_out(cbx_1__1__70_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__70_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__70_ccff_tail)
  );


  cbx_1__1_
  cbx_8__11_
  (
    .clk_1_S_out(clk_1_wires[167]),
    .clk_1_N_out(clk_1_wires[166]),
    .clk_1_W_in(clk_1_wires[162]),
    .prog_clk_1_S_out(prog_clk_1_wires[167]),
    .prog_clk_1_N_out(prog_clk_1_wires[166]),
    .prog_clk_1_W_in(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[324]),
    .config_enable_S_out(config_enableWires[582]),
    .config_enable_E_out(config_enableWires[581]),
    .config_enable_W_in(config_enableWires[580]),
    .sc_head_N_out(sc_headWires[206]),
    .sc_head_S_in(sc_headWires[205]),
    .pReset_S_out(pResetWires[582]),
    .pReset_E_out(pResetWires[581]),
    .pReset_W_in(pResetWires[580]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[87]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[87]),
    .chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__48_ccff_tail),
    .chanx_left_out(cbx_1__1__71_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__71_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__71_ccff_tail)
  );


  cbx_1__1_
  cbx_9__1_
  (
    .clk_1_S_out(clk_1_wires[172]),
    .clk_1_N_out(clk_1_wires[171]),
    .clk_1_E_in(clk_1_wires[170]),
    .prog_clk_1_S_out(prog_clk_1_wires[172]),
    .prog_clk_1_N_out(prog_clk_1_wires[171]),
    .prog_clk_1_E_in(prog_clk_1_wires[170]),
    .prog_clk_0_N_in(prog_clk_0_wires[332]),
    .config_enable_S_out(config_enableWires[96]),
    .config_enable_E_out(config_enableWires[95]),
    .config_enable_W_in(config_enableWires[94]),
    .sc_head_S_out(sc_headWires[232]),
    .sc_head_N_in(sc_headWires[231]),
    .pReset_S_out(pResetWires[96]),
    .pReset_E_out(pResetWires[95]),
    .pReset_W_in(pResetWires[94]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[88]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[88]),
    .chanx_left_in(sb_1__1__49_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__49_ccff_tail),
    .chanx_left_out(cbx_1__1__72_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__72_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__72_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__72_ccff_tail)
  );


  cbx_1__1_
  cbx_9__2_
  (
    .clk_2_E_out(clk_2_wires[70]),
    .clk_2_W_in(clk_2_wires[69]),
    .prog_clk_2_E_out(prog_clk_2_wires[70]),
    .prog_clk_2_W_in(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[335]),
    .config_enable_S_out(config_enableWires[145]),
    .config_enable_E_out(config_enableWires[144]),
    .config_enable_W_in(config_enableWires[143]),
    .sc_head_S_out(sc_headWires[230]),
    .sc_head_N_in(sc_headWires[229]),
    .pReset_S_out(pResetWires[145]),
    .pReset_E_out(pResetWires[144]),
    .pReset_W_in(pResetWires[143]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[89]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[89]),
    .chanx_left_in(sb_2__2__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__8_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__6_ccff_tail),
    .chanx_left_out(cbx_1__1__73_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__73_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__73_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__73_ccff_tail)
  );


  cbx_1__1_
  cbx_9__4_
  (
    .clk_2_E_out(clk_2_wires[79]),
    .clk_2_W_in(clk_2_wires[78]),
    .prog_clk_2_E_out(prog_clk_2_wires[79]),
    .prog_clk_2_W_in(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[341]),
    .config_enable_S_out(config_enableWires[243]),
    .config_enable_E_out(config_enableWires[242]),
    .config_enable_W_in(config_enableWires[241]),
    .sc_head_S_out(sc_headWires[226]),
    .sc_head_N_in(sc_headWires[225]),
    .pReset_S_out(pResetWires[243]),
    .pReset_E_out(pResetWires[242]),
    .pReset_W_in(pResetWires[241]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[91]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[91]),
    .chanx_left_in(sb_1__1__50_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__50_ccff_tail),
    .chanx_left_out(cbx_1__1__74_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__74_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__74_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__74_ccff_tail)
  );


  cbx_1__1_
  cbx_9__5_
  (
    .clk_1_S_out(clk_1_wires[186]),
    .clk_1_N_out(clk_1_wires[185]),
    .clk_1_E_in(clk_1_wires[184]),
    .prog_clk_1_S_out(prog_clk_1_wires[186]),
    .prog_clk_1_N_out(prog_clk_1_wires[185]),
    .prog_clk_1_E_in(prog_clk_1_wires[184]),
    .prog_clk_0_N_in(prog_clk_0_wires[344]),
    .config_enable_S_out(config_enableWires[292]),
    .config_enable_E_out(config_enableWires[291]),
    .config_enable_W_in(config_enableWires[290]),
    .sc_head_S_out(sc_headWires[224]),
    .sc_head_N_in(sc_headWires[223]),
    .pReset_S_out(pResetWires[292]),
    .pReset_E_out(pResetWires[291]),
    .pReset_W_in(pResetWires[290]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[92]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[92]),
    .chanx_left_in(sb_1__1__51_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__51_ccff_tail),
    .chanx_left_out(cbx_1__1__75_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__75_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__75_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__75_ccff_tail)
  );


  cbx_1__1_
  cbx_9__6_
  (
    .clk_3_E_out(clk_3_wires[45]),
    .clk_3_W_in(clk_3_wires[44]),
    .prog_clk_3_E_out(prog_clk_3_wires[45]),
    .prog_clk_3_W_in(prog_clk_3_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[347]),
    .config_enable_S_out(config_enableWires[341]),
    .config_enable_E_out(config_enableWires[340]),
    .config_enable_W_in(config_enableWires[339]),
    .sc_head_S_out(sc_headWires[222]),
    .sc_head_N_in(sc_headWires[221]),
    .pReset_S_out(pResetWires[341]),
    .pReset_E_out(pResetWires[340]),
    .pReset_W_in(pResetWires[339]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[93]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[93]),
    .chanx_left_in(sb_1__1__52_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__52_ccff_tail),
    .chanx_left_out(cbx_1__1__76_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__76_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__76_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__76_ccff_tail)
  );


  cbx_1__1_
  cbx_9__7_
  (
    .clk_1_S_out(clk_1_wires[193]),
    .clk_1_N_out(clk_1_wires[192]),
    .clk_1_E_in(clk_1_wires[191]),
    .prog_clk_1_S_out(prog_clk_1_wires[193]),
    .prog_clk_1_N_out(prog_clk_1_wires[192]),
    .prog_clk_1_E_in(prog_clk_1_wires[191]),
    .prog_clk_0_N_in(prog_clk_0_wires[350]),
    .config_enable_S_out(config_enableWires[390]),
    .config_enable_E_out(config_enableWires[389]),
    .config_enable_W_in(config_enableWires[388]),
    .sc_head_S_out(sc_headWires[220]),
    .sc_head_N_in(sc_headWires[219]),
    .pReset_S_out(pResetWires[390]),
    .pReset_E_out(pResetWires[389]),
    .pReset_W_in(pResetWires[388]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[94]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[94]),
    .chanx_left_in(sb_1__1__53_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__53_ccff_tail),
    .chanx_left_out(cbx_1__1__77_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__77_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__77_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__77_ccff_tail)
  );


  cbx_1__1_
  cbx_9__8_
  (
    .clk_2_E_out(clk_2_wires[92]),
    .clk_2_W_in(clk_2_wires[91]),
    .prog_clk_2_E_out(prog_clk_2_wires[92]),
    .prog_clk_2_W_in(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[353]),
    .config_enable_S_out(config_enableWires[439]),
    .config_enable_E_out(config_enableWires[438]),
    .config_enable_W_in(config_enableWires[437]),
    .sc_head_S_out(sc_headWires[218]),
    .sc_head_N_in(sc_headWires[217]),
    .pReset_S_out(pResetWires[439]),
    .pReset_E_out(pResetWires[438]),
    .pReset_W_in(pResetWires[437]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[95]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[95]),
    .chanx_left_in(sb_1__1__54_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__54_ccff_tail),
    .chanx_left_out(cbx_1__1__78_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__78_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__78_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__78_ccff_tail)
  );


  cbx_1__1_
  cbx_9__9_
  (
    .clk_1_S_out(clk_1_wires[200]),
    .clk_1_N_out(clk_1_wires[199]),
    .clk_1_E_in(clk_1_wires[198]),
    .prog_clk_1_S_out(prog_clk_1_wires[200]),
    .prog_clk_1_N_out(prog_clk_1_wires[199]),
    .prog_clk_1_E_in(prog_clk_1_wires[198]),
    .prog_clk_0_N_in(prog_clk_0_wires[356]),
    .config_enable_S_out(config_enableWires[488]),
    .config_enable_E_out(config_enableWires[487]),
    .config_enable_W_in(config_enableWires[486]),
    .sc_head_S_out(sc_headWires[216]),
    .sc_head_N_in(sc_headWires[215]),
    .pReset_S_out(pResetWires[488]),
    .pReset_E_out(pResetWires[487]),
    .pReset_W_in(pResetWires[486]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[96]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[96]),
    .chanx_left_in(sb_2__2__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__9_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__7_ccff_tail),
    .chanx_left_out(cbx_1__1__79_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__79_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__79_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__79_ccff_tail)
  );


  cbx_1__1_
  cbx_9__11_
  (
    .clk_1_S_out(clk_1_wires[207]),
    .clk_1_N_out(clk_1_wires[206]),
    .clk_1_E_in(clk_1_wires[205]),
    .prog_clk_1_S_out(prog_clk_1_wires[207]),
    .prog_clk_1_N_out(prog_clk_1_wires[206]),
    .prog_clk_1_E_in(prog_clk_1_wires[205]),
    .prog_clk_0_N_in(prog_clk_0_wires[362]),
    .config_enable_S_out(config_enableWires[586]),
    .config_enable_E_out(config_enableWires[585]),
    .config_enable_W_in(config_enableWires[584]),
    .sc_head_S_out(sc_headWires[212]),
    .sc_head_N_in(sc_headWires[211]),
    .pReset_S_out(pResetWires[586]),
    .pReset_E_out(pResetWires[585]),
    .pReset_W_in(pResetWires[584]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[98]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[98]),
    .chanx_left_in(sb_1__1__55_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__55_ccff_tail),
    .chanx_left_out(cbx_1__1__80_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__80_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__80_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__80_ccff_tail)
  );


  cbx_1__1_
  cbx_10__1_
  (
    .clk_1_S_out(clk_1_wires[174]),
    .clk_1_N_out(clk_1_wires[173]),
    .clk_1_W_in(clk_1_wires[169]),
    .prog_clk_1_S_out(prog_clk_1_wires[174]),
    .prog_clk_1_N_out(prog_clk_1_wires[173]),
    .prog_clk_1_W_in(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[370]),
    .config_enable_S_out(config_enableWires[100]),
    .config_enable_E_out(config_enableWires[99]),
    .config_enable_W_in(config_enableWires[98]),
    .sc_head_N_out(sc_headWires[238]),
    .sc_head_S_in(sc_headWires[237]),
    .pReset_S_out(pResetWires[100]),
    .pReset_E_out(pResetWires[99]),
    .pReset_W_in(pResetWires[98]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[99]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[99]),
    .chanx_left_in(sb_1__1__56_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__56_ccff_tail),
    .chanx_left_out(cbx_1__1__81_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__81_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__81_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__81_ccff_tail)
  );


  cbx_1__1_
  cbx_10__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[373]),
    .config_enable_S_out(config_enableWires[149]),
    .config_enable_E_out(config_enableWires[148]),
    .config_enable_W_in(config_enableWires[147]),
    .sc_head_N_out(sc_headWires[240]),
    .sc_head_S_in(sc_headWires[239]),
    .pReset_S_out(pResetWires[149]),
    .pReset_E_out(pResetWires[148]),
    .pReset_W_in(pResetWires[147]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[100]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[100]),
    .chanx_left_in(sb_1__2__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__8_ccff_tail),
    .chanx_left_out(cbx_1__1__82_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__82_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__82_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__82_ccff_tail)
  );


  cbx_1__1_
  cbx_10__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[379]),
    .config_enable_S_out(config_enableWires[247]),
    .config_enable_E_out(config_enableWires[246]),
    .config_enable_W_in(config_enableWires[245]),
    .sc_head_N_out(sc_headWires[244]),
    .sc_head_S_in(sc_headWires[243]),
    .pReset_S_out(pResetWires[247]),
    .pReset_E_out(pResetWires[246]),
    .pReset_W_in(pResetWires[245]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[102]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[102]),
    .chanx_left_in(sb_1__1__57_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__57_ccff_tail),
    .chanx_left_out(cbx_1__1__83_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__83_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__83_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__83_ccff_tail)
  );


  cbx_1__1_
  cbx_10__5_
  (
    .clk_1_S_out(clk_1_wires[188]),
    .clk_1_N_out(clk_1_wires[187]),
    .clk_1_W_in(clk_1_wires[183]),
    .prog_clk_1_S_out(prog_clk_1_wires[188]),
    .prog_clk_1_N_out(prog_clk_1_wires[187]),
    .prog_clk_1_W_in(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[382]),
    .config_enable_S_out(config_enableWires[296]),
    .config_enable_E_out(config_enableWires[295]),
    .config_enable_W_in(config_enableWires[294]),
    .sc_head_N_out(sc_headWires[246]),
    .sc_head_S_in(sc_headWires[245]),
    .pReset_S_out(pResetWires[296]),
    .pReset_E_out(pResetWires[295]),
    .pReset_W_in(pResetWires[294]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[103]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[103]),
    .chanx_left_in(sb_1__1__58_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__58_ccff_tail),
    .chanx_left_out(cbx_1__1__84_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__84_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__84_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__84_ccff_tail)
  );


  cbx_1__1_
  cbx_10__6_
  (
    .clk_3_E_out(clk_3_wires[49]),
    .clk_3_W_in(clk_3_wires[48]),
    .prog_clk_3_E_out(prog_clk_3_wires[49]),
    .prog_clk_3_W_in(prog_clk_3_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[385]),
    .config_enable_S_out(config_enableWires[345]),
    .config_enable_E_out(config_enableWires[344]),
    .config_enable_W_in(config_enableWires[343]),
    .sc_head_N_out(sc_headWires[248]),
    .sc_head_S_in(sc_headWires[247]),
    .pReset_S_out(pResetWires[345]),
    .pReset_E_out(pResetWires[344]),
    .pReset_W_in(pResetWires[343]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[104]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[104]),
    .chanx_left_in(sb_1__1__59_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__59_ccff_tail),
    .chanx_left_out(cbx_1__1__85_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__85_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__85_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__85_ccff_tail)
  );


  cbx_1__1_
  cbx_10__7_
  (
    .clk_1_S_out(clk_1_wires[195]),
    .clk_1_N_out(clk_1_wires[194]),
    .clk_1_W_in(clk_1_wires[190]),
    .prog_clk_1_S_out(prog_clk_1_wires[195]),
    .prog_clk_1_N_out(prog_clk_1_wires[194]),
    .prog_clk_1_W_in(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[388]),
    .config_enable_S_out(config_enableWires[394]),
    .config_enable_E_out(config_enableWires[393]),
    .config_enable_W_in(config_enableWires[392]),
    .sc_head_N_out(sc_headWires[250]),
    .sc_head_S_in(sc_headWires[249]),
    .pReset_S_out(pResetWires[394]),
    .pReset_E_out(pResetWires[393]),
    .pReset_W_in(pResetWires[392]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[105]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[105]),
    .chanx_left_in(sb_1__1__60_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__60_ccff_tail),
    .chanx_left_out(cbx_1__1__86_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__86_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__86_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__86_ccff_tail)
  );


  cbx_1__1_
  cbx_10__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[391]),
    .config_enable_S_out(config_enableWires[443]),
    .config_enable_E_out(config_enableWires[442]),
    .config_enable_W_in(config_enableWires[441]),
    .sc_head_N_out(sc_headWires[252]),
    .sc_head_S_in(sc_headWires[251]),
    .pReset_S_out(pResetWires[443]),
    .pReset_E_out(pResetWires[442]),
    .pReset_W_in(pResetWires[441]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[106]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[106]),
    .chanx_left_in(sb_1__1__61_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__61_ccff_tail),
    .chanx_left_out(cbx_1__1__87_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__87_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__87_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__87_ccff_tail)
  );


  cbx_1__1_
  cbx_10__9_
  (
    .clk_1_S_out(clk_1_wires[202]),
    .clk_1_N_out(clk_1_wires[201]),
    .clk_1_W_in(clk_1_wires[197]),
    .prog_clk_1_S_out(prog_clk_1_wires[202]),
    .prog_clk_1_N_out(prog_clk_1_wires[201]),
    .prog_clk_1_W_in(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[394]),
    .config_enable_S_out(config_enableWires[492]),
    .config_enable_E_out(config_enableWires[491]),
    .config_enable_W_in(config_enableWires[490]),
    .sc_head_N_out(sc_headWires[254]),
    .sc_head_S_in(sc_headWires[253]),
    .pReset_S_out(pResetWires[492]),
    .pReset_E_out(pResetWires[491]),
    .pReset_W_in(pResetWires[490]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[107]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[107]),
    .chanx_left_in(sb_1__2__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__2__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__9_ccff_tail),
    .chanx_left_out(cbx_1__1__88_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__88_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__88_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__88_ccff_tail)
  );


  cbx_1__1_
  cbx_10__11_
  (
    .clk_1_S_out(clk_1_wires[209]),
    .clk_1_N_out(clk_1_wires[208]),
    .clk_1_W_in(clk_1_wires[204]),
    .prog_clk_1_S_out(prog_clk_1_wires[209]),
    .prog_clk_1_N_out(prog_clk_1_wires[208]),
    .prog_clk_1_W_in(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[400]),
    .config_enable_S_out(config_enableWires[590]),
    .config_enable_E_out(config_enableWires[589]),
    .config_enable_W_in(config_enableWires[588]),
    .sc_head_N_out(sc_headWires[258]),
    .sc_head_S_in(sc_headWires[257]),
    .pReset_S_out(pResetWires[590]),
    .pReset_E_out(pResetWires[589]),
    .pReset_W_in(pResetWires[588]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[109]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[109]),
    .chanx_left_in(sb_1__1__62_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__62_ccff_tail),
    .chanx_left_out(cbx_1__1__89_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__89_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__89_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__89_ccff_tail)
  );


  cbx_1__1_
  cbx_11__1_
  (
    .clk_1_S_out(clk_1_wires[214]),
    .clk_1_N_out(clk_1_wires[213]),
    .clk_1_E_in(clk_1_wires[212]),
    .prog_clk_1_S_out(prog_clk_1_wires[214]),
    .prog_clk_1_N_out(prog_clk_1_wires[213]),
    .prog_clk_1_E_in(prog_clk_1_wires[212]),
    .prog_clk_0_N_in(prog_clk_0_wires[408]),
    .config_enable_S_out(config_enableWires[104]),
    .config_enable_E_out(config_enableWires[103]),
    .config_enable_W_in(config_enableWires[102]),
    .sc_head_S_out(sc_headWires[284]),
    .sc_head_N_in(sc_headWires[283]),
    .pReset_S_out(pResetWires[104]),
    .pReset_E_out(pResetWires[103]),
    .pReset_W_in(pResetWires[102]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[110]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[110]),
    .chanx_left_in(sb_1__1__63_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__63_ccff_tail),
    .chanx_left_out(cbx_1__1__90_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__90_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__90_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__90_ccff_tail)
  );


  cbx_1__1_
  cbx_11__2_
  (
    .clk_2_W_in(clk_2_wires[114]),
    .clk_2_E_out(clk_2_wires[113]),
    .prog_clk_2_W_in(prog_clk_2_wires[114]),
    .prog_clk_2_E_out(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[411]),
    .config_enable_S_out(config_enableWires[153]),
    .config_enable_E_out(config_enableWires[152]),
    .config_enable_W_in(config_enableWires[151]),
    .sc_head_S_out(sc_headWires[282]),
    .sc_head_N_in(sc_headWires[281]),
    .pReset_S_out(pResetWires[153]),
    .pReset_E_out(pResetWires[152]),
    .pReset_W_in(pResetWires[151]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[111]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[111]),
    .chanx_left_in(sb_2__2__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__10_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__8_ccff_tail),
    .chanx_left_out(cbx_1__1__91_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__91_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__91_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__91_ccff_tail)
  );


  cbx_1__1_
  cbx_11__4_
  (
    .clk_2_W_in(clk_2_wires[119]),
    .clk_2_E_out(clk_2_wires[118]),
    .prog_clk_2_W_in(prog_clk_2_wires[119]),
    .prog_clk_2_E_out(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[417]),
    .config_enable_S_out(config_enableWires[251]),
    .config_enable_E_out(config_enableWires[250]),
    .config_enable_W_in(config_enableWires[249]),
    .sc_head_S_out(sc_headWires[278]),
    .sc_head_N_in(sc_headWires[277]),
    .pReset_S_out(pResetWires[251]),
    .pReset_E_out(pResetWires[250]),
    .pReset_W_in(pResetWires[249]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[113]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[113]),
    .chanx_left_in(sb_1__1__64_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__64_ccff_tail),
    .chanx_left_out(cbx_1__1__92_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__92_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__92_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__92_ccff_tail)
  );


  cbx_1__1_
  cbx_11__5_
  (
    .clk_1_S_out(clk_1_wires[228]),
    .clk_1_N_out(clk_1_wires[227]),
    .clk_1_E_in(clk_1_wires[226]),
    .prog_clk_1_S_out(prog_clk_1_wires[228]),
    .prog_clk_1_N_out(prog_clk_1_wires[227]),
    .prog_clk_1_E_in(prog_clk_1_wires[226]),
    .prog_clk_0_N_in(prog_clk_0_wires[420]),
    .config_enable_S_out(config_enableWires[300]),
    .config_enable_E_out(config_enableWires[299]),
    .config_enable_W_in(config_enableWires[298]),
    .sc_head_S_out(sc_headWires[276]),
    .sc_head_N_in(sc_headWires[275]),
    .pReset_S_out(pResetWires[300]),
    .pReset_E_out(pResetWires[299]),
    .pReset_W_in(pResetWires[298]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[114]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[114]),
    .chanx_left_in(sb_1__1__65_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__65_ccff_tail),
    .chanx_left_out(cbx_1__1__93_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__93_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__93_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__93_ccff_tail)
  );


  cbx_1__1_
  cbx_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[423]),
    .config_enable_S_out(config_enableWires[349]),
    .config_enable_E_out(config_enableWires[348]),
    .config_enable_W_in(config_enableWires[347]),
    .sc_head_S_out(sc_headWires[274]),
    .sc_head_N_in(sc_headWires[273]),
    .pReset_S_out(pResetWires[349]),
    .pReset_E_out(pResetWires[348]),
    .pReset_W_in(pResetWires[347]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[115]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[115]),
    .chanx_left_in(sb_1__1__66_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__66_ccff_tail),
    .chanx_left_out(cbx_1__1__94_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__94_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__94_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__94_ccff_tail)
  );


  cbx_1__1_
  cbx_11__7_
  (
    .clk_1_S_out(clk_1_wires[235]),
    .clk_1_N_out(clk_1_wires[234]),
    .clk_1_E_in(clk_1_wires[233]),
    .prog_clk_1_S_out(prog_clk_1_wires[235]),
    .prog_clk_1_N_out(prog_clk_1_wires[234]),
    .prog_clk_1_E_in(prog_clk_1_wires[233]),
    .prog_clk_0_N_in(prog_clk_0_wires[426]),
    .config_enable_S_out(config_enableWires[398]),
    .config_enable_E_out(config_enableWires[397]),
    .config_enable_W_in(config_enableWires[396]),
    .sc_head_S_out(sc_headWires[272]),
    .sc_head_N_in(sc_headWires[271]),
    .pReset_S_out(pResetWires[398]),
    .pReset_E_out(pResetWires[397]),
    .pReset_W_in(pResetWires[396]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[116]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[116]),
    .chanx_left_in(sb_1__1__67_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__67_ccff_tail),
    .chanx_left_out(cbx_1__1__95_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__95_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__95_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__95_ccff_tail)
  );


  cbx_1__1_
  cbx_11__8_
  (
    .clk_2_W_in(clk_2_wires[126]),
    .clk_2_E_out(clk_2_wires[125]),
    .prog_clk_2_W_in(prog_clk_2_wires[126]),
    .prog_clk_2_E_out(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[429]),
    .config_enable_S_out(config_enableWires[447]),
    .config_enable_E_out(config_enableWires[446]),
    .config_enable_W_in(config_enableWires[445]),
    .sc_head_S_out(sc_headWires[270]),
    .sc_head_N_in(sc_headWires[269]),
    .pReset_S_out(pResetWires[447]),
    .pReset_E_out(pResetWires[446]),
    .pReset_W_in(pResetWires[445]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[117]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[117]),
    .chanx_left_in(sb_1__1__68_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__68_ccff_tail),
    .chanx_left_out(cbx_1__1__96_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__96_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__96_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__96_ccff_tail)
  );


  cbx_1__1_
  cbx_11__9_
  (
    .clk_1_S_out(clk_1_wires[242]),
    .clk_1_N_out(clk_1_wires[241]),
    .clk_1_E_in(clk_1_wires[240]),
    .prog_clk_1_S_out(prog_clk_1_wires[242]),
    .prog_clk_1_N_out(prog_clk_1_wires[241]),
    .prog_clk_1_E_in(prog_clk_1_wires[240]),
    .prog_clk_0_N_in(prog_clk_0_wires[432]),
    .config_enable_S_out(config_enableWires[496]),
    .config_enable_E_out(config_enableWires[495]),
    .config_enable_W_in(config_enableWires[494]),
    .sc_head_S_out(sc_headWires[268]),
    .sc_head_N_in(sc_headWires[267]),
    .pReset_S_out(pResetWires[496]),
    .pReset_E_out(pResetWires[495]),
    .pReset_W_in(pResetWires[494]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[118]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[118]),
    .chanx_left_in(sb_2__2__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__2__11_chanx_left_out[0:19]),
    .ccff_head(sb_2__2__9_ccff_tail),
    .chanx_left_out(cbx_1__1__97_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__97_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__97_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__97_ccff_tail)
  );


  cbx_1__1_
  cbx_11__11_
  (
    .clk_1_S_out(clk_1_wires[249]),
    .clk_1_N_out(clk_1_wires[248]),
    .clk_1_E_in(clk_1_wires[247]),
    .prog_clk_1_S_out(prog_clk_1_wires[249]),
    .prog_clk_1_N_out(prog_clk_1_wires[248]),
    .prog_clk_1_E_in(prog_clk_1_wires[247]),
    .prog_clk_0_N_in(prog_clk_0_wires[438]),
    .config_enable_S_out(config_enableWires[594]),
    .config_enable_E_out(config_enableWires[593]),
    .config_enable_W_in(config_enableWires[592]),
    .sc_head_S_out(sc_headWires[264]),
    .sc_head_N_in(sc_headWires[263]),
    .pReset_S_out(pResetWires[594]),
    .pReset_E_out(pResetWires[593]),
    .pReset_W_in(pResetWires[592]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[120]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[120]),
    .chanx_left_in(sb_1__1__69_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__69_ccff_tail),
    .chanx_left_out(cbx_1__1__98_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__98_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__98_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__98_ccff_tail)
  );


  cbx_1__1_
  cbx_12__1_
  (
    .clk_1_S_out(clk_1_wires[216]),
    .clk_1_N_out(clk_1_wires[215]),
    .clk_1_W_in(clk_1_wires[211]),
    .prog_clk_1_S_out(prog_clk_1_wires[216]),
    .prog_clk_1_N_out(prog_clk_1_wires[215]),
    .prog_clk_1_W_in(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[446]),
    .config_enable_S_out(config_enableWires[108]),
    .config_enable_E_out(config_enableWires[107]),
    .config_enable_W_in(config_enableWires[106]),
    .sc_head_N_out(sc_headWires[290]),
    .sc_head_S_in(sc_headWires[289]),
    .pReset_S_out(pResetWires[108]),
    .pReset_E_out(pResetWires[107]),
    .pReset_W_in(pResetWires[106]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[121]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[121]),
    .chanx_left_in(sb_1__1__70_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__70_ccff_tail),
    .chanx_left_out(cbx_1__1__99_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__99_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__99_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__99_ccff_tail)
  );


  cbx_1__1_
  cbx_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[449]),
    .config_enable_S_out(config_enableWires[157]),
    .config_enable_E_out(config_enableWires[156]),
    .config_enable_W_in(config_enableWires[155]),
    .sc_head_N_out(sc_headWires[292]),
    .sc_head_S_in(sc_headWires[291]),
    .pReset_S_out(pResetWires[157]),
    .pReset_E_out(pResetWires[156]),
    .pReset_W_in(pResetWires[155]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[122]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[122]),
    .chanx_left_in(sb_1__2__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__2__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__10_ccff_tail),
    .chanx_left_out(cbx_1__1__100_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__100_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__100_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__100_ccff_tail)
  );


  cbx_1__1_
  cbx_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[455]),
    .config_enable_S_out(config_enableWires[255]),
    .config_enable_E_out(config_enableWires[254]),
    .config_enable_W_in(config_enableWires[253]),
    .sc_head_N_out(sc_headWires[296]),
    .sc_head_S_in(sc_headWires[295]),
    .pReset_S_out(pResetWires[255]),
    .pReset_E_out(pResetWires[254]),
    .pReset_W_in(pResetWires[253]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[124]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[124]),
    .chanx_left_in(sb_1__1__71_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__71_ccff_tail),
    .chanx_left_out(cbx_1__1__101_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__101_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__101_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__101_ccff_tail)
  );


  cbx_1__1_
  cbx_12__5_
  (
    .clk_1_S_out(clk_1_wires[230]),
    .clk_1_N_out(clk_1_wires[229]),
    .clk_1_W_in(clk_1_wires[225]),
    .prog_clk_1_S_out(prog_clk_1_wires[230]),
    .prog_clk_1_N_out(prog_clk_1_wires[229]),
    .prog_clk_1_W_in(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[458]),
    .config_enable_S_out(config_enableWires[304]),
    .config_enable_E_out(config_enableWires[303]),
    .config_enable_W_in(config_enableWires[302]),
    .sc_head_N_out(sc_headWires[298]),
    .sc_head_S_in(sc_headWires[297]),
    .pReset_S_out(pResetWires[304]),
    .pReset_E_out(pResetWires[303]),
    .pReset_W_in(pResetWires[302]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[125]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[125]),
    .chanx_left_in(sb_1__1__72_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__72_ccff_tail),
    .chanx_left_out(cbx_1__1__102_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__102_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__102_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__102_ccff_tail)
  );


  cbx_1__1_
  cbx_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[461]),
    .config_enable_S_out(config_enableWires[353]),
    .config_enable_E_out(config_enableWires[352]),
    .config_enable_W_in(config_enableWires[351]),
    .sc_head_N_out(sc_headWires[300]),
    .sc_head_S_in(sc_headWires[299]),
    .pReset_S_out(pResetWires[353]),
    .pReset_E_out(pResetWires[352]),
    .pReset_W_in(pResetWires[351]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[126]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[126]),
    .chanx_left_in(sb_1__1__73_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__73_ccff_tail),
    .chanx_left_out(cbx_1__1__103_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__103_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__103_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__103_ccff_tail)
  );


  cbx_1__1_
  cbx_12__7_
  (
    .clk_1_S_out(clk_1_wires[237]),
    .clk_1_N_out(clk_1_wires[236]),
    .clk_1_W_in(clk_1_wires[232]),
    .prog_clk_1_S_out(prog_clk_1_wires[237]),
    .prog_clk_1_N_out(prog_clk_1_wires[236]),
    .prog_clk_1_W_in(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[464]),
    .config_enable_S_out(config_enableWires[402]),
    .config_enable_E_out(config_enableWires[401]),
    .config_enable_W_in(config_enableWires[400]),
    .sc_head_N_out(sc_headWires[302]),
    .sc_head_S_in(sc_headWires[301]),
    .pReset_S_out(pResetWires[402]),
    .pReset_E_out(pResetWires[401]),
    .pReset_W_in(pResetWires[400]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[127]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[127]),
    .chanx_left_in(sb_1__1__74_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__74_ccff_tail),
    .chanx_left_out(cbx_1__1__104_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__104_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__104_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__104_ccff_tail)
  );


  cbx_1__1_
  cbx_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[467]),
    .config_enable_S_out(config_enableWires[451]),
    .config_enable_E_out(config_enableWires[450]),
    .config_enable_W_in(config_enableWires[449]),
    .sc_head_N_out(sc_headWires[304]),
    .sc_head_S_in(sc_headWires[303]),
    .pReset_S_out(pResetWires[451]),
    .pReset_E_out(pResetWires[450]),
    .pReset_W_in(pResetWires[449]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[128]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[128]),
    .chanx_left_in(sb_1__1__75_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__75_ccff_tail),
    .chanx_left_out(cbx_1__1__105_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__105_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__105_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__105_ccff_tail)
  );


  cbx_1__1_
  cbx_12__9_
  (
    .clk_1_S_out(clk_1_wires[244]),
    .clk_1_N_out(clk_1_wires[243]),
    .clk_1_W_in(clk_1_wires[239]),
    .prog_clk_1_S_out(prog_clk_1_wires[244]),
    .prog_clk_1_N_out(prog_clk_1_wires[243]),
    .prog_clk_1_W_in(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[470]),
    .config_enable_S_out(config_enableWires[500]),
    .config_enable_E_out(config_enableWires[499]),
    .config_enable_W_in(config_enableWires[498]),
    .sc_head_N_out(sc_headWires[306]),
    .sc_head_S_in(sc_headWires[305]),
    .pReset_S_out(pResetWires[500]),
    .pReset_E_out(pResetWires[499]),
    .pReset_W_in(pResetWires[498]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[129]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[129]),
    .chanx_left_in(sb_1__2__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__2__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__2__11_ccff_tail),
    .chanx_left_out(cbx_1__1__106_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__106_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__106_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__106_ccff_tail)
  );


  cbx_1__1_
  cbx_12__11_
  (
    .clk_1_S_out(clk_1_wires[251]),
    .clk_1_N_out(clk_1_wires[250]),
    .clk_1_W_in(clk_1_wires[246]),
    .prog_clk_1_S_out(prog_clk_1_wires[251]),
    .prog_clk_1_N_out(prog_clk_1_wires[250]),
    .prog_clk_1_W_in(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[476]),
    .config_enable_S_out(config_enableWires[598]),
    .config_enable_E_out(config_enableWires[597]),
    .config_enable_W_in(config_enableWires[596]),
    .sc_head_N_out(sc_headWires[310]),
    .sc_head_S_in(sc_headWires[309]),
    .pReset_S_out(pResetWires[598]),
    .pReset_E_out(pResetWires[597]),
    .pReset_W_in(pResetWires[596]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[131]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[131]),
    .chanx_left_in(sb_1__1__76_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__76_ccff_tail),
    .chanx_left_out(cbx_1__1__107_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__107_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_6_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_7_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__107_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
    .ccff_tail(cbx_1__1__107_ccff_tail)
  );


  cbx_1__3_
  cbx_1__3_
  (
    .clk_1_S_out(clk_1_wires[11]),
    .clk_1_N_out(clk_1_wires[10]),
    .clk_1_E_in(clk_1_wires[9]),
    .prog_clk_1_S_out(prog_clk_1_wires[11]),
    .prog_clk_1_N_out(prog_clk_1_wires[10]),
    .prog_clk_1_E_in(prog_clk_1_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[16]),
    .prog_clk_0_W_out(prog_clk_0_wires[15]),
    .config_enable_S_out(config_enableWires[161]),
    .config_enable_E_in(config_enableWires[160]),
    .config_enable_W_out(config_enableWires[159]),
    .sc_head_S_out(sc_headWires[20]),
    .sc_head_N_in(sc_headWires[19]),
    .pReset_S_out(pResetWires[161]),
    .pReset_E_in(pResetWires[160]),
    .pReset_W_out(pResetWires[159]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[2]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[2]),
    .chanx_left_in(sb_0__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_0__3__0_ccff_tail),
    .chanx_left_out(cbx_1__3__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__0_ccff_tail)
  );


  cbx_1__3_
  cbx_1__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[51]),
    .prog_clk_0_W_out(prog_clk_0_wires[50]),
    .config_enable_S_out(config_enableWires[504]),
    .config_enable_E_in(config_enableWires[503]),
    .config_enable_W_out(config_enableWires[502]),
    .sc_head_S_out(sc_headWires[6]),
    .sc_head_N_in(sc_headWires[5]),
    .pReset_S_out(pResetWires[504]),
    .pReset_E_in(pResetWires[503]),
    .pReset_W_out(pResetWires[502]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[9]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[9]),
    .chanx_left_in(sb_0__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_0__3__1_ccff_tail),
    .chanx_left_out(cbx_1__3__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__1_ccff_tail)
  );


  cbx_1__3_
  cbx_3__3_
  (
    .clk_1_S_out(clk_1_wires[53]),
    .clk_1_N_out(clk_1_wires[52]),
    .clk_1_E_in(clk_1_wires[51]),
    .prog_clk_1_S_out(prog_clk_1_wires[53]),
    .prog_clk_1_N_out(prog_clk_1_wires[52]),
    .prog_clk_1_E_in(prog_clk_1_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[110]),
    .config_enable_S_out(config_enableWires[170]),
    .config_enable_E_in(config_enableWires[169]),
    .config_enable_W_out(config_enableWires[168]),
    .sc_head_S_out(sc_headWires[72]),
    .sc_head_N_in(sc_headWires[71]),
    .pReset_S_out(pResetWires[170]),
    .pReset_E_in(pResetWires[169]),
    .pReset_W_out(pResetWires[168]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[24]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[24]),
    .chanx_left_in(sb_2__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__2_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__0_ccff_tail),
    .chanx_left_out(cbx_1__3__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__2_ccff_tail)
  );


  cbx_1__3_
  cbx_3__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[131]),
    .config_enable_S_out(config_enableWires[513]),
    .config_enable_E_in(config_enableWires[512]),
    .config_enable_W_out(config_enableWires[511]),
    .sc_head_S_out(sc_headWires[58]),
    .sc_head_N_in(sc_headWires[57]),
    .pReset_S_out(pResetWires[513]),
    .pReset_E_in(pResetWires[512]),
    .pReset_W_out(pResetWires[511]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[31]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[31]),
    .chanx_left_in(sb_2__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__3_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__1_ccff_tail),
    .chanx_left_out(cbx_1__3__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__3_ccff_tail)
  );


  cbx_1__3_
  cbx_5__3_
  (
    .clk_1_S_out(clk_1_wires[95]),
    .clk_1_N_out(clk_1_wires[94]),
    .clk_1_E_in(clk_1_wires[93]),
    .prog_clk_1_S_out(prog_clk_1_wires[95]),
    .prog_clk_1_N_out(prog_clk_1_wires[94]),
    .prog_clk_1_E_in(prog_clk_1_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[186]),
    .config_enable_S_out(config_enableWires[178]),
    .config_enable_E_in(config_enableWires[177]),
    .config_enable_W_out(config_enableWires[176]),
    .sc_head_S_out(sc_headWires[124]),
    .sc_head_N_in(sc_headWires[123]),
    .pReset_S_out(pResetWires[178]),
    .pReset_E_in(pResetWires[177]),
    .pReset_W_out(pResetWires[176]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[46]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[46]),
    .chanx_left_in(sb_2__3__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__4_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__2_ccff_tail),
    .chanx_left_out(cbx_1__3__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__4_ccff_tail)
  );


  cbx_1__3_
  cbx_5__10_
  (
    .clk_2_E_out(clk_2_wires[61]),
    .clk_2_W_in(clk_2_wires[60]),
    .prog_clk_2_E_out(prog_clk_2_wires[61]),
    .prog_clk_2_W_in(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[207]),
    .config_enable_S_out(config_enableWires[521]),
    .config_enable_E_in(config_enableWires[520]),
    .config_enable_W_out(config_enableWires[519]),
    .sc_head_S_out(sc_headWires[110]),
    .sc_head_N_in(sc_headWires[109]),
    .pReset_S_out(pResetWires[521]),
    .pReset_E_in(pResetWires[520]),
    .pReset_W_out(pResetWires[519]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[53]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[53]),
    .chanx_left_in(sb_2__3__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__5_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__3_ccff_tail),
    .chanx_left_out(cbx_1__3__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__5_ccff_tail)
  );


  cbx_1__3_
  cbx_7__3_
  (
    .clk_1_S_out(clk_1_wires[137]),
    .clk_1_N_out(clk_1_wires[136]),
    .clk_1_E_in(clk_1_wires[135]),
    .prog_clk_1_S_out(prog_clk_1_wires[137]),
    .prog_clk_1_N_out(prog_clk_1_wires[136]),
    .prog_clk_1_E_in(prog_clk_1_wires[135]),
    .prog_clk_0_N_in(prog_clk_0_wires[262]),
    .config_enable_S_out(config_enableWires[186]),
    .config_enable_E_out(config_enableWires[185]),
    .config_enable_W_in(config_enableWires[184]),
    .sc_head_S_out(sc_headWires[176]),
    .sc_head_N_in(sc_headWires[175]),
    .pReset_S_out(pResetWires[186]),
    .pReset_E_out(pResetWires[185]),
    .pReset_W_in(pResetWires[184]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[68]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[68]),
    .chanx_left_in(sb_2__3__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__6_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__4_ccff_tail),
    .chanx_left_out(cbx_1__3__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__6_ccff_tail)
  );


  cbx_1__3_
  cbx_7__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[283]),
    .config_enable_S_out(config_enableWires[529]),
    .config_enable_E_out(config_enableWires[528]),
    .config_enable_W_in(config_enableWires[527]),
    .sc_head_S_out(sc_headWires[162]),
    .sc_head_N_in(sc_headWires[161]),
    .pReset_S_out(pResetWires[529]),
    .pReset_E_out(pResetWires[528]),
    .pReset_W_in(pResetWires[527]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[75]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[75]),
    .chanx_left_in(sb_2__3__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__7_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__5_ccff_tail),
    .chanx_left_out(cbx_1__3__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__7_ccff_tail)
  );


  cbx_1__3_
  cbx_9__3_
  (
    .clk_1_S_out(clk_1_wires[179]),
    .clk_1_N_out(clk_1_wires[178]),
    .clk_1_E_in(clk_1_wires[177]),
    .prog_clk_1_S_out(prog_clk_1_wires[179]),
    .prog_clk_1_N_out(prog_clk_1_wires[178]),
    .prog_clk_1_E_in(prog_clk_1_wires[177]),
    .prog_clk_0_N_in(prog_clk_0_wires[338]),
    .config_enable_S_out(config_enableWires[194]),
    .config_enable_E_out(config_enableWires[193]),
    .config_enable_W_in(config_enableWires[192]),
    .sc_head_S_out(sc_headWires[228]),
    .sc_head_N_in(sc_headWires[227]),
    .pReset_S_out(pResetWires[194]),
    .pReset_E_out(pResetWires[193]),
    .pReset_W_in(pResetWires[192]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[90]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[90]),
    .chanx_left_in(sb_2__3__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__8_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__6_ccff_tail),
    .chanx_left_out(cbx_1__3__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__8_ccff_tail)
  );


  cbx_1__3_
  cbx_9__10_
  (
    .clk_2_E_out(clk_2_wires[105]),
    .clk_2_W_in(clk_2_wires[104]),
    .prog_clk_2_E_out(prog_clk_2_wires[105]),
    .prog_clk_2_W_in(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[359]),
    .config_enable_S_out(config_enableWires[537]),
    .config_enable_E_out(config_enableWires[536]),
    .config_enable_W_in(config_enableWires[535]),
    .sc_head_S_out(sc_headWires[214]),
    .sc_head_N_in(sc_headWires[213]),
    .pReset_S_out(pResetWires[537]),
    .pReset_E_out(pResetWires[536]),
    .pReset_W_in(pResetWires[535]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[97]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[97]),
    .chanx_left_in(sb_2__3__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__9_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__7_ccff_tail),
    .chanx_left_out(cbx_1__3__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__9_ccff_tail)
  );


  cbx_1__3_
  cbx_11__3_
  (
    .clk_1_S_out(clk_1_wires[221]),
    .clk_1_N_out(clk_1_wires[220]),
    .clk_1_E_in(clk_1_wires[219]),
    .prog_clk_1_S_out(prog_clk_1_wires[221]),
    .prog_clk_1_N_out(prog_clk_1_wires[220]),
    .prog_clk_1_E_in(prog_clk_1_wires[219]),
    .prog_clk_0_N_in(prog_clk_0_wires[414]),
    .config_enable_S_out(config_enableWires[202]),
    .config_enable_E_out(config_enableWires[201]),
    .config_enable_W_in(config_enableWires[200]),
    .sc_head_S_out(sc_headWires[280]),
    .sc_head_N_in(sc_headWires[279]),
    .pReset_S_out(pResetWires[202]),
    .pReset_E_out(pResetWires[201]),
    .pReset_W_in(pResetWires[200]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[112]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[112]),
    .chanx_left_in(sb_2__3__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__10_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__8_ccff_tail),
    .chanx_left_out(cbx_1__3__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__10_ccff_tail)
  );


  cbx_1__3_
  cbx_11__10_
  (
    .clk_2_W_in(clk_2_wires[133]),
    .clk_2_E_out(clk_2_wires[132]),
    .prog_clk_2_W_in(prog_clk_2_wires[133]),
    .prog_clk_2_E_out(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[435]),
    .config_enable_S_out(config_enableWires[545]),
    .config_enable_E_out(config_enableWires[544]),
    .config_enable_W_in(config_enableWires[543]),
    .sc_head_S_out(sc_headWires[266]),
    .sc_head_N_in(sc_headWires[265]),
    .pReset_S_out(pResetWires[545]),
    .pReset_E_out(pResetWires[544]),
    .pReset_W_in(pResetWires[543]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[119]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[119]),
    .chanx_left_in(sb_2__3__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__3__11_chanx_left_out[0:19]),
    .ccff_head(sb_2__3__9_ccff_tail),
    .chanx_left_out(cbx_1__3__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__3__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
    .bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
    .ccff_tail(cbx_1__3__11_ccff_tail)
  );


  cbx_1__4_
  cbx_1__12_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[62]),
    .prog_clk_0_S_in(prog_clk_0_wires[59]),
    .config_enable_S_out(config_enableWires[602]),
    .config_enable_E_in(config_enableWires[601]),
    .config_enable_W_out(config_enableWires[600]),
    .sc_head_S_out(sc_headWires[2]),
    .sc_head_W_in(sc_headWires[1]),
    .pReset_S_out(pResetWires[602]),
    .pReset_E_in(pResetWires[601]),
    .pReset_W_out(pResetWires[600]),
    .chanx_left_in(sb_0__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_head(grid_clb_9_ccff_tail),
    .chanx_left_out(cbx_1__12__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__0_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[0]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[0]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[0]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_0_ccff_tail)
  );


  cbx_1__4_
  cbx_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[99]),
    .config_enable_S_out(config_enableWires[606]),
    .config_enable_E_in(config_enableWires[605]),
    .config_enable_W_out(config_enableWires[604]),
    .sc_head_E_out(sc_headWires[52]),
    .sc_head_S_in(sc_headWires[51]),
    .pReset_S_out(pResetWires[606]),
    .pReset_E_in(pResetWires[605]),
    .pReset_W_out(pResetWires[604]),
    .chanx_left_in(sb_1__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_head(grid_clb_19_ccff_tail),
    .chanx_left_out(cbx_1__12__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__1_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[1]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[1]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[1]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_1_ccff_tail)
  );


  cbx_1__4_
  cbx_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[137]),
    .config_enable_S_out(config_enableWires[609]),
    .config_enable_E_in(config_enableWires[608]),
    .config_enable_W_out(config_enableWires[607]),
    .sc_head_S_out(sc_headWires[54]),
    .sc_head_W_in(sc_headWires[53]),
    .pReset_S_out(pResetWires[609]),
    .pReset_E_in(pResetWires[608]),
    .pReset_W_out(pResetWires[607]),
    .chanx_left_in(sb_1__12__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_head(grid_clb_29_ccff_tail),
    .chanx_left_out(cbx_1__12__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__2_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[2]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[2]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[2]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_2_ccff_tail)
  );


  cbx_1__4_
  cbx_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[175]),
    .config_enable_S_out(config_enableWires[612]),
    .config_enable_E_in(config_enableWires[611]),
    .config_enable_W_out(config_enableWires[610]),
    .sc_head_E_out(sc_headWires[104]),
    .sc_head_S_in(sc_headWires[103]),
    .pReset_S_out(pResetWires[612]),
    .pReset_E_in(pResetWires[611]),
    .pReset_W_out(pResetWires[610]),
    .chanx_left_in(sb_1__12__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_head(grid_clb_39_ccff_tail),
    .chanx_left_out(cbx_1__12__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__3_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[3]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[3]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[3]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_3_ccff_tail)
  );


  cbx_1__4_
  cbx_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[213]),
    .config_enable_S_out(config_enableWires[615]),
    .config_enable_E_in(config_enableWires[614]),
    .config_enable_W_out(config_enableWires[613]),
    .sc_head_S_out(sc_headWires[106]),
    .sc_head_W_in(sc_headWires[105]),
    .pReset_S_out(pResetWires[615]),
    .pReset_E_in(pResetWires[614]),
    .pReset_W_out(pResetWires[613]),
    .chanx_left_in(sb_1__12__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_head(grid_clb_49_ccff_tail),
    .chanx_left_out(cbx_1__12__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__4_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[4]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[4]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[4]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_4_ccff_tail)
  );


  cbx_1__4_
  cbx_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[251]),
    .config_enable_S_out(config_enableWires[618]),
    .config_enable_E_in(config_enableWires[617]),
    .config_enable_W_out(config_enableWires[616]),
    .sc_head_E_out(sc_headWires[156]),
    .sc_head_S_in(sc_headWires[155]),
    .pReset_S_out(pResetWires[618]),
    .pReset_E_in(pResetWires[617]),
    .pReset_W_out(pResetWires[616]),
    .chanx_left_in(sb_1__12__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_head(grid_clb_59_ccff_tail),
    .chanx_left_out(cbx_1__12__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__5_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[5]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[5]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[5]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_5_ccff_tail)
  );


  cbx_1__4_
  cbx_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[289]),
    .config_enable_S_out(config_enableWires[621]),
    .config_enable_E_out(config_enableWires[620]),
    .config_enable_W_in(config_enableWires[619]),
    .sc_head_S_out(sc_headWires[158]),
    .sc_head_W_in(sc_headWires[157]),
    .pReset_S_out(pResetWires[621]),
    .pReset_E_out(pResetWires[620]),
    .pReset_W_in(pResetWires[619]),
    .chanx_left_in(sb_1__12__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_head(grid_clb_69_ccff_tail),
    .chanx_left_out(cbx_1__12__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__6_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[6]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[6]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[6]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_6_ccff_tail)
  );


  cbx_1__4_
  cbx_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[327]),
    .config_enable_S_out(config_enableWires[624]),
    .config_enable_E_out(config_enableWires[623]),
    .config_enable_W_in(config_enableWires[622]),
    .sc_head_E_out(sc_headWires[208]),
    .sc_head_S_in(sc_headWires[207]),
    .pReset_S_out(pResetWires[624]),
    .pReset_E_out(pResetWires[623]),
    .pReset_W_in(pResetWires[622]),
    .chanx_left_in(sb_1__12__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_head(grid_clb_79_ccff_tail),
    .chanx_left_out(cbx_1__12__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__7_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[7]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[7]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[7]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_7_ccff_tail)
  );


  cbx_1__4_
  cbx_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[365]),
    .config_enable_S_out(config_enableWires[627]),
    .config_enable_E_out(config_enableWires[626]),
    .config_enable_W_in(config_enableWires[625]),
    .sc_head_S_out(sc_headWires[210]),
    .sc_head_W_in(sc_headWires[209]),
    .pReset_S_out(pResetWires[627]),
    .pReset_E_out(pResetWires[626]),
    .pReset_W_in(pResetWires[625]),
    .chanx_left_in(sb_1__12__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_head(grid_clb_89_ccff_tail),
    .chanx_left_out(cbx_1__12__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__8_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[8]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[8]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[8]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_8_ccff_tail)
  );


  cbx_1__4_
  cbx_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[403]),
    .config_enable_S_out(config_enableWires[630]),
    .config_enable_E_out(config_enableWires[629]),
    .config_enable_W_in(config_enableWires[628]),
    .sc_head_E_out(sc_headWires[260]),
    .sc_head_S_in(sc_headWires[259]),
    .pReset_S_out(pResetWires[630]),
    .pReset_E_out(pResetWires[629]),
    .pReset_W_in(pResetWires[628]),
    .chanx_left_in(sb_1__12__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_head(grid_clb_99_ccff_tail),
    .chanx_left_out(cbx_1__12__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__9_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[9]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[9]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[9]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_9_ccff_tail)
  );


  cbx_1__4_
  cbx_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[441]),
    .config_enable_S_out(config_enableWires[633]),
    .config_enable_E_out(config_enableWires[632]),
    .config_enable_W_in(config_enableWires[631]),
    .sc_head_S_out(sc_headWires[262]),
    .sc_head_W_in(sc_headWires[261]),
    .pReset_S_out(pResetWires[633]),
    .pReset_E_out(pResetWires[632]),
    .pReset_W_in(pResetWires[631]),
    .chanx_left_in(sb_1__12__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_head(grid_clb_109_ccff_tail),
    .chanx_left_out(cbx_1__12__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__10_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[10]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[10]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[10]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_10_ccff_tail)
  );


  cbx_1__4_
  cbx_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[479]),
    .config_enable_S_out(config_enableWires[636]),
    .config_enable_E_out(config_enableWires[635]),
    .config_enable_W_in(config_enableWires[634]),
    .sc_head_E_out(sc_headWires[312]),
    .sc_head_S_in(sc_headWires[311]),
    .pReset_S_out(pResetWires[636]),
    .pReset_E_out(pResetWires[635]),
    .pReset_W_in(pResetWires[634]),
    .chanx_left_in(sb_1__12__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_head(grid_clb_119_ccff_tail),
    .chanx_left_out(cbx_1__12__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__11_chanx_right_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[11]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[11]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[11]),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_top_top_11_ccff_tail)
  );


  cbx_2__3_
  cbx_2__3_
  (
    .clk_1_S_out(clk_1_wires[13]),
    .clk_1_N_out(clk_1_wires[12]),
    .clk_1_W_in(clk_1_wires[8]),
    .prog_clk_1_S_out(prog_clk_1_wires[13]),
    .prog_clk_1_N_out(prog_clk_1_wires[12]),
    .prog_clk_1_W_in(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[72]),
    .config_enable_S_out(config_enableWires[166]),
    .config_enable_E_in(config_enableWires[165]),
    .config_enable_W_out(config_enableWires[164]),
    .sc_head_N_out(sc_headWires[34]),
    .sc_head_S_in(sc_headWires[33]),
    .pReset_S_out(pResetWires[166]),
    .pReset_E_in(pResetWires[165]),
    .pReset_W_out(pResetWires[164]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[13]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[13]),
    .chanx_left_in(sb_1__3__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__0_ccff_tail),
    .chanx_left_out(cbx_2__3__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__0_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__0_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__0_ccff_tail)
  );


  cbx_2__3_
  cbx_2__10_
  (
    .clk_2_E_in(clk_2_wires[21]),
    .clk_2_W_out(clk_2_wires[20]),
    .prog_clk_2_E_in(prog_clk_2_wires[21]),
    .prog_clk_2_W_out(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[93]),
    .config_enable_S_out(config_enableWires[509]),
    .config_enable_E_in(config_enableWires[508]),
    .config_enable_W_out(config_enableWires[507]),
    .sc_head_N_out(sc_headWires[48]),
    .sc_head_S_in(sc_headWires[47]),
    .pReset_S_out(pResetWires[509]),
    .pReset_E_in(pResetWires[508]),
    .pReset_W_out(pResetWires[507]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[20]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[20]),
    .chanx_left_in(sb_1__3__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__1_ccff_tail),
    .chanx_left_out(cbx_2__3__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__1_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__1_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__1_ccff_tail)
  );


  cbx_2__3_
  cbx_4__3_
  (
    .clk_1_S_out(clk_1_wires[55]),
    .clk_1_N_out(clk_1_wires[54]),
    .clk_1_W_in(clk_1_wires[50]),
    .prog_clk_1_S_out(prog_clk_1_wires[55]),
    .prog_clk_1_N_out(prog_clk_1_wires[54]),
    .prog_clk_1_W_in(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[148]),
    .config_enable_S_out(config_enableWires[174]),
    .config_enable_E_in(config_enableWires[173]),
    .config_enable_W_out(config_enableWires[172]),
    .sc_head_N_out(sc_headWires[86]),
    .sc_head_S_in(sc_headWires[85]),
    .pReset_S_out(pResetWires[174]),
    .pReset_E_in(pResetWires[173]),
    .pReset_W_out(pResetWires[172]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[35]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[35]),
    .chanx_left_in(sb_1__3__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__2_ccff_tail),
    .chanx_left_out(cbx_2__3__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__2_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__2_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__2_ccff_tail)
  );


  cbx_2__3_
  cbx_4__10_
  (
    .clk_2_W_out(clk_2_wires[63]),
    .clk_2_E_in(clk_2_wires[62]),
    .prog_clk_2_W_out(prog_clk_2_wires[63]),
    .prog_clk_2_E_in(prog_clk_2_wires[62]),
    .prog_clk_0_N_in(prog_clk_0_wires[169]),
    .config_enable_S_out(config_enableWires[517]),
    .config_enable_E_in(config_enableWires[516]),
    .config_enable_W_out(config_enableWires[515]),
    .sc_head_N_out(sc_headWires[100]),
    .sc_head_S_in(sc_headWires[99]),
    .pReset_S_out(pResetWires[517]),
    .pReset_E_in(pResetWires[516]),
    .pReset_W_out(pResetWires[515]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[42]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[42]),
    .chanx_left_in(sb_1__3__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__3_ccff_tail),
    .chanx_left_out(cbx_2__3__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__3_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__3_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__3_ccff_tail)
  );


  cbx_2__3_
  cbx_6__3_
  (
    .clk_1_S_out(clk_1_wires[97]),
    .clk_1_N_out(clk_1_wires[96]),
    .clk_1_W_in(clk_1_wires[92]),
    .prog_clk_1_S_out(prog_clk_1_wires[97]),
    .prog_clk_1_N_out(prog_clk_1_wires[96]),
    .prog_clk_1_W_in(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[224]),
    .config_enable_S_out(config_enableWires[182]),
    .config_enable_E_in(config_enableWires[181]),
    .config_enable_W_out(config_enableWires[180]),
    .sc_head_N_out(sc_headWires[138]),
    .sc_head_S_in(sc_headWires[137]),
    .pReset_S_out(pResetWires[182]),
    .pReset_E_in(pResetWires[181]),
    .pReset_W_out(pResetWires[180]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[57]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[57]),
    .chanx_left_in(sb_1__3__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__4_ccff_tail),
    .chanx_left_out(cbx_2__3__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__4_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__4_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__4_ccff_tail)
  );


  cbx_2__3_
  cbx_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[245]),
    .config_enable_S_out(config_enableWires[525]),
    .config_enable_E_in(config_enableWires[524]),
    .config_enable_W_out(config_enableWires[523]),
    .sc_head_N_out(sc_headWires[152]),
    .sc_head_S_in(sc_headWires[151]),
    .pReset_S_out(pResetWires[525]),
    .pReset_E_in(pResetWires[524]),
    .pReset_W_out(pResetWires[523]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[64]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[64]),
    .chanx_left_in(sb_1__3__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__5_ccff_tail),
    .chanx_left_out(cbx_2__3__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__5_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__5_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__5_ccff_tail)
  );


  cbx_2__3_
  cbx_8__3_
  (
    .clk_1_S_out(clk_1_wires[139]),
    .clk_1_N_out(clk_1_wires[138]),
    .clk_1_W_in(clk_1_wires[134]),
    .prog_clk_1_S_out(prog_clk_1_wires[139]),
    .prog_clk_1_N_out(prog_clk_1_wires[138]),
    .prog_clk_1_W_in(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[300]),
    .config_enable_S_out(config_enableWires[190]),
    .config_enable_E_out(config_enableWires[189]),
    .config_enable_W_in(config_enableWires[188]),
    .sc_head_N_out(sc_headWires[190]),
    .sc_head_S_in(sc_headWires[189]),
    .pReset_S_out(pResetWires[190]),
    .pReset_E_out(pResetWires[189]),
    .pReset_W_in(pResetWires[188]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[79]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[79]),
    .chanx_left_in(sb_1__3__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__6_ccff_tail),
    .chanx_left_out(cbx_2__3__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__6_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__6_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__6_ccff_tail)
  );


  cbx_2__3_
  cbx_8__10_
  (
    .clk_2_W_out(clk_2_wires[107]),
    .clk_2_E_in(clk_2_wires[106]),
    .prog_clk_2_W_out(prog_clk_2_wires[107]),
    .prog_clk_2_E_in(prog_clk_2_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[321]),
    .config_enable_S_out(config_enableWires[533]),
    .config_enable_E_out(config_enableWires[532]),
    .config_enable_W_in(config_enableWires[531]),
    .sc_head_N_out(sc_headWires[204]),
    .sc_head_S_in(sc_headWires[203]),
    .pReset_S_out(pResetWires[533]),
    .pReset_E_out(pResetWires[532]),
    .pReset_W_in(pResetWires[531]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[86]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[86]),
    .chanx_left_in(sb_1__3__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__7_ccff_tail),
    .chanx_left_out(cbx_2__3__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__7_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__7_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__7_ccff_tail)
  );


  cbx_2__3_
  cbx_10__3_
  (
    .clk_1_S_out(clk_1_wires[181]),
    .clk_1_N_out(clk_1_wires[180]),
    .clk_1_W_in(clk_1_wires[176]),
    .prog_clk_1_S_out(prog_clk_1_wires[181]),
    .prog_clk_1_N_out(prog_clk_1_wires[180]),
    .prog_clk_1_W_in(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[376]),
    .config_enable_S_out(config_enableWires[198]),
    .config_enable_E_out(config_enableWires[197]),
    .config_enable_W_in(config_enableWires[196]),
    .sc_head_N_out(sc_headWires[242]),
    .sc_head_S_in(sc_headWires[241]),
    .pReset_S_out(pResetWires[198]),
    .pReset_E_out(pResetWires[197]),
    .pReset_W_in(pResetWires[196]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[101]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[101]),
    .chanx_left_in(sb_1__3__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__8_ccff_tail),
    .chanx_left_out(cbx_2__3__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__8_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__8_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__8_ccff_tail)
  );


  cbx_2__3_
  cbx_10__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[397]),
    .config_enable_S_out(config_enableWires[541]),
    .config_enable_E_out(config_enableWires[540]),
    .config_enable_W_in(config_enableWires[539]),
    .sc_head_N_out(sc_headWires[256]),
    .sc_head_S_in(sc_headWires[255]),
    .pReset_S_out(pResetWires[541]),
    .pReset_E_out(pResetWires[540]),
    .pReset_W_in(pResetWires[539]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[108]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[108]),
    .chanx_left_in(sb_1__3__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_2__3__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__9_ccff_tail),
    .chanx_left_out(cbx_2__3__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__9_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__9_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__9_ccff_tail)
  );


  cbx_2__3_
  cbx_12__3_
  (
    .clk_1_S_out(clk_1_wires[223]),
    .clk_1_N_out(clk_1_wires[222]),
    .clk_1_W_in(clk_1_wires[218]),
    .prog_clk_1_S_out(prog_clk_1_wires[223]),
    .prog_clk_1_N_out(prog_clk_1_wires[222]),
    .prog_clk_1_W_in(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[452]),
    .config_enable_S_out(config_enableWires[206]),
    .config_enable_E_out(config_enableWires[205]),
    .config_enable_W_in(config_enableWires[204]),
    .sc_head_N_out(sc_headWires[294]),
    .sc_head_S_in(sc_headWires[293]),
    .pReset_S_out(pResetWires[206]),
    .pReset_E_out(pResetWires[205]),
    .pReset_W_in(pResetWires[204]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[123]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[123]),
    .chanx_left_in(sb_1__3__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__3__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__10_ccff_tail),
    .chanx_left_out(cbx_2__3__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__10_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__10_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__10_ccff_tail)
  );


  cbx_2__3_
  cbx_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[473]),
    .config_enable_S_out(config_enableWires[549]),
    .config_enable_E_out(config_enableWires[548]),
    .config_enable_W_in(config_enableWires[547]),
    .sc_head_N_out(sc_headWires[308]),
    .sc_head_S_in(sc_headWires[307]),
    .pReset_S_out(pResetWires[549]),
    .pReset_E_out(pResetWires[548]),
    .pReset_W_in(pResetWires[547]),
    .REG_OUT_FEEDTHROUGH(reg_out__feedthrough_wires[130]),
    .REG_IN_FEEDTHROUGH(reg_in_feedthrough_wires[130]),
    .chanx_left_in(sb_1__3__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__3__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__3__11_ccff_tail),
    .chanx_left_out(cbx_2__3__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_2__3__11_chanx_right_out[0:19]),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_a_11_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_6_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_7_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_8_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_9_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_10_),
    .bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_(cbx_2__3__11_bottom_grid_top_width_1_height_0_subtile_0__pin_b_11_),
    .ccff_tail(cbx_2__3__11_ccff_tail)
  );


  cby_0__1_
  cby_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[3]),
    .config_enable_N_in(config_enableWires[64]),
    .pReset_N_in(pResetWires[64]),
    .chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_0_ccff_tail),
    .chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__0_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[132]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[132]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[132]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_0_ccff_tail)
  );


  cby_0__1_
  cby_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[9]),
    .config_enable_N_in(config_enableWires[113]),
    .pReset_N_in(pResetWires[113]),
    .chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_1_ccff_tail),
    .chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__1_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[133]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[133]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[133]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_1_ccff_tail)
  );


  cby_0__1_
  cby_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[14]),
    .config_enable_N_in(config_enableWires[162]),
    .pReset_N_in(pResetWires[162]),
    .chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__3__0_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_0_ccff_tail),
    .chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__2_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[134]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[134]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[134]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_2_ccff_tail)
  );


  cby_0__1_
  cby_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[19]),
    .config_enable_N_in(config_enableWires[211]),
    .pReset_N_in(pResetWires[211]),
    .chany_bottom_in(sb_0__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_2_ccff_tail),
    .chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__3_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[135]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[135]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[135]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_3_ccff_tail)
  );


  cby_0__1_
  cby_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[24]),
    .config_enable_N_in(config_enableWires[260]),
    .pReset_N_in(pResetWires[260]),
    .chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_3_ccff_tail),
    .chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__4_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[136]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[136]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[136]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_4_ccff_tail)
  );


  cby_0__1_
  cby_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[29]),
    .config_enable_N_in(config_enableWires[309]),
    .pReset_N_in(pResetWires[309]),
    .chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_4_ccff_tail),
    .chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__5_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[137]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[137]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[137]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_5_ccff_tail)
  );


  cby_0__1_
  cby_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[34]),
    .config_enable_N_in(config_enableWires[358]),
    .pReset_N_in(pResetWires[358]),
    .chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_5_ccff_tail),
    .chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__6_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[138]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[138]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[138]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_6_ccff_tail)
  );


  cby_0__1_
  cby_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[39]),
    .config_enable_N_in(config_enableWires[407]),
    .pReset_N_in(pResetWires[407]),
    .chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_6_ccff_tail),
    .chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__7_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[139]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[139]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[139]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_7_ccff_tail)
  );


  cby_0__1_
  cby_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[44]),
    .config_enable_N_in(config_enableWires[456]),
    .pReset_N_in(pResetWires[456]),
    .chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_7_ccff_tail),
    .chany_bottom_out(cby_0__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__8_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[140]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[140]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[140]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_8_ccff_tail)
  );


  cby_0__1_
  cby_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[49]),
    .config_enable_N_in(config_enableWires[505]),
    .pReset_N_in(pResetWires[505]),
    .chany_bottom_in(sb_0__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_0__3__1_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_1_ccff_tail),
    .chany_bottom_out(cby_0__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__9_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[141]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[141]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[141]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_9_ccff_tail)
  );


  cby_0__1_
  cby_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[54]),
    .config_enable_N_in(config_enableWires[554]),
    .pReset_N_in(pResetWires[554]),
    .chany_bottom_in(sb_0__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_8_ccff_tail),
    .chany_bottom_out(cby_0__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__10_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[142]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[142]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[142]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_10_ccff_tail)
  );


  cby_0__1_
  cby_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[61]),
    .config_enable_N_in(config_enableWires[603]),
    .pReset_N_in(pResetWires[603]),
    .chany_bottom_in(sb_0__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__12__0_ccff_tail),
    .chany_bottom_out(cby_0__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__11_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[143]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[143]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[143]),
    .right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_left_left_11_ccff_tail)
  );


  cby_1__1_
  cby_1__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[2]),
    .prog_clk_0_W_in(prog_clk_0_wires[1]),
    .config_enable_S_in(config_enableWires[27]),
    .reset_E_in(resetWires[26]),
    .reset_W_out(resetWires[24]),
    .Test_en_E_in(Test_enWires[26]),
    .Test_en_W_out(Test_enWires[24]),
    .pReset_S_in(pResetWires[27]),
    .chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_10_ccff_tail),
    .chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__0_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__0_ccff_tail)
  );


  cby_1__1_
  cby_1__2_
  (
    .clk_2_S_out(clk_2_wires[4]),
    .clk_2_N_in(clk_2_wires[3]),
    .prog_clk_2_S_out(prog_clk_2_wires[4]),
    .prog_clk_2_N_in(prog_clk_2_wires[3]),
    .prog_clk_0_S_out(prog_clk_0_wires[8]),
    .prog_clk_0_W_in(prog_clk_0_wires[7]),
    .config_enable_S_in(config_enableWires[65]),
    .reset_E_in(resetWires[48]),
    .reset_W_out(resetWires[46]),
    .Test_en_E_in(Test_enWires[48]),
    .Test_en_W_out(Test_enWires[46]),
    .pReset_S_in(pResetWires[65]),
    .chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_11_ccff_tail),
    .chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__1_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__1_ccff_tail)
  );


  cby_1__1_
  cby_1__4_
  (
    .clk_2_S_out(clk_2_wires[11]),
    .clk_2_N_in(clk_2_wires[10]),
    .prog_clk_2_S_out(prog_clk_2_wires[11]),
    .prog_clk_2_N_in(prog_clk_2_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[18]),
    .prog_clk_0_W_in(prog_clk_0_wires[17]),
    .config_enable_S_in(config_enableWires[163]),
    .reset_E_in(resetWires[92]),
    .reset_W_out(resetWires[90]),
    .Test_en_E_in(Test_enWires[92]),
    .Test_en_W_out(Test_enWires[90]),
    .pReset_S_in(pResetWires[163]),
    .chany_bottom_in(sb_1__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_12_ccff_tail),
    .chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__2_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__2_ccff_tail)
  );


  cby_1__1_
  cby_1__5_
  (
    .clk_2_N_out(clk_2_wires[9]),
    .clk_2_S_in(clk_2_wires[8]),
    .prog_clk_2_N_out(prog_clk_2_wires[9]),
    .prog_clk_2_S_in(prog_clk_2_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[23]),
    .prog_clk_0_W_in(prog_clk_0_wires[22]),
    .config_enable_S_in(config_enableWires[212]),
    .reset_E_in(resetWires[114]),
    .reset_W_out(resetWires[112]),
    .Test_en_E_in(Test_enWires[114]),
    .Test_en_W_out(Test_enWires[112]),
    .pReset_S_in(pResetWires[212]),
    .chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_13_ccff_tail),
    .chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__3_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__3_ccff_tail)
  );


  cby_1__1_
  cby_1__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[28]),
    .prog_clk_0_W_in(prog_clk_0_wires[27]),
    .config_enable_S_in(config_enableWires[261]),
    .reset_E_in(resetWires[136]),
    .reset_W_out(resetWires[134]),
    .Test_en_E_in(Test_enWires[136]),
    .Test_en_W_out(Test_enWires[134]),
    .pReset_S_in(pResetWires[261]),
    .chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_14_ccff_tail),
    .chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__4_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__4_ccff_tail)
  );


  cby_1__1_
  cby_1__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[33]),
    .prog_clk_0_W_in(prog_clk_0_wires[32]),
    .config_enable_S_in(config_enableWires[310]),
    .reset_E_in(resetWires[158]),
    .reset_W_out(resetWires[156]),
    .Test_en_E_in(Test_enWires[158]),
    .Test_en_W_out(Test_enWires[156]),
    .pReset_S_in(pResetWires[310]),
    .chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_15_ccff_tail),
    .chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__5_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__5_ccff_tail)
  );


  cby_1__1_
  cby_1__8_
  (
    .clk_2_S_out(clk_2_wires[18]),
    .clk_2_N_in(clk_2_wires[17]),
    .prog_clk_2_S_out(prog_clk_2_wires[18]),
    .prog_clk_2_N_in(prog_clk_2_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[38]),
    .prog_clk_0_W_in(prog_clk_0_wires[37]),
    .config_enable_S_in(config_enableWires[359]),
    .reset_E_in(resetWires[180]),
    .reset_W_out(resetWires[178]),
    .Test_en_E_in(Test_enWires[180]),
    .Test_en_W_out(Test_enWires[178]),
    .pReset_S_in(pResetWires[359]),
    .chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_16_ccff_tail),
    .chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__6_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__6_ccff_tail)
  );


  cby_1__1_
  cby_1__9_
  (
    .clk_2_N_out(clk_2_wires[16]),
    .clk_2_S_in(clk_2_wires[15]),
    .prog_clk_2_N_out(prog_clk_2_wires[16]),
    .prog_clk_2_S_in(prog_clk_2_wires[15]),
    .prog_clk_0_S_out(prog_clk_0_wires[43]),
    .prog_clk_0_W_in(prog_clk_0_wires[42]),
    .config_enable_S_in(config_enableWires[408]),
    .reset_E_in(resetWires[202]),
    .reset_W_out(resetWires[200]),
    .Test_en_E_in(Test_enWires[202]),
    .Test_en_W_out(Test_enWires[200]),
    .pReset_S_in(pResetWires[408]),
    .chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_17_ccff_tail),
    .chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__7_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__7_ccff_tail)
  );


  cby_1__1_
  cby_1__11_
  (
    .clk_2_N_out(clk_2_wires[23]),
    .clk_2_S_in(clk_2_wires[22]),
    .prog_clk_2_N_out(prog_clk_2_wires[23]),
    .prog_clk_2_S_in(prog_clk_2_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[53]),
    .prog_clk_0_W_in(prog_clk_0_wires[52]),
    .config_enable_S_in(config_enableWires[506]),
    .reset_E_in(resetWires[246]),
    .reset_W_out(resetWires[244]),
    .Test_en_E_in(Test_enWires[246]),
    .Test_en_W_out(Test_enWires[244]),
    .pReset_S_in(pResetWires[506]),
    .chany_bottom_in(sb_1__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_18_ccff_tail),
    .chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__8_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__8_ccff_tail)
  );


  cby_1__1_
  cby_1__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[60]),
    .prog_clk_0_S_out(prog_clk_0_wires[58]),
    .prog_clk_0_W_in(prog_clk_0_wires[57]),
    .config_enable_S_in(config_enableWires[555]),
    .reset_E_in(resetWires[268]),
    .reset_W_out(resetWires[266]),
    .Test_en_E_in(Test_enWires[268]),
    .Test_en_W_out(Test_enWires[266]),
    .pReset_S_in(pResetWires[555]),
    .chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__0_ccff_tail),
    .chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__9_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__9_ccff_tail)
  );


  cby_1__1_
  cby_2__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[65]),
    .prog_clk_0_W_in(prog_clk_0_wires[64]),
    .config_enable_S_in(config_enableWires[30]),
    .reset_E_in(resetWires[28]),
    .reset_W_out(resetWires[25]),
    .Test_en_E_in(Test_enWires[28]),
    .Test_en_W_out(Test_enWires[25]),
    .pReset_S_in(pResetWires[30]),
    .chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_20_ccff_tail),
    .chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__10_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__10_ccff_tail)
  );


  cby_1__1_
  cby_2__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[68]),
    .prog_clk_0_W_in(prog_clk_0_wires[67]),
    .config_enable_S_in(config_enableWires[69]),
    .reset_E_in(resetWires[50]),
    .reset_W_out(resetWires[47]),
    .Test_en_E_in(Test_enWires[50]),
    .Test_en_W_out(Test_enWires[47]),
    .pReset_S_in(pResetWires[69]),
    .chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_21_ccff_tail),
    .chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__11_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__11_ccff_tail)
  );


  cby_1__1_
  cby_2__4_
  (
    .clk_3_S_out(clk_3_wires[65]),
    .clk_3_N_in(clk_3_wires[64]),
    .prog_clk_3_S_out(prog_clk_3_wires[65]),
    .prog_clk_3_N_in(prog_clk_3_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[74]),
    .prog_clk_0_W_in(prog_clk_0_wires[73]),
    .config_enable_S_in(config_enableWires[167]),
    .reset_E_in(resetWires[94]),
    .reset_W_out(resetWires[91]),
    .Test_en_E_in(Test_enWires[94]),
    .Test_en_W_out(Test_enWires[91]),
    .pReset_S_in(pResetWires[167]),
    .chany_bottom_in(sb_2__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_22_ccff_tail),
    .chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__12_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__12_ccff_tail)
  );


  cby_1__1_
  cby_2__5_
  (
    .clk_3_S_out(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[58]),
    .prog_clk_3_S_out(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[58]),
    .prog_clk_0_S_out(prog_clk_0_wires[77]),
    .prog_clk_0_W_in(prog_clk_0_wires[76]),
    .config_enable_S_in(config_enableWires[216]),
    .reset_E_in(resetWires[116]),
    .reset_W_out(resetWires[113]),
    .Test_en_E_in(Test_enWires[116]),
    .Test_en_W_out(Test_enWires[113]),
    .pReset_S_in(pResetWires[216]),
    .chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_23_ccff_tail),
    .chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__13_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__13_ccff_tail)
  );


  cby_1__1_
  cby_2__6_
  (
    .clk_3_S_out(clk_3_wires[55]),
    .clk_3_N_in(clk_3_wires[54]),
    .prog_clk_3_S_out(prog_clk_3_wires[55]),
    .prog_clk_3_N_in(prog_clk_3_wires[54]),
    .prog_clk_0_S_out(prog_clk_0_wires[80]),
    .prog_clk_0_W_in(prog_clk_0_wires[79]),
    .config_enable_S_in(config_enableWires[265]),
    .reset_E_in(resetWires[138]),
    .reset_W_out(resetWires[135]),
    .Test_en_E_in(Test_enWires[138]),
    .Test_en_W_out(Test_enWires[135]),
    .pReset_S_in(pResetWires[265]),
    .chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_24_ccff_tail),
    .chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__14_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__14_ccff_tail)
  );


  cby_1__1_
  cby_2__7_
  (
    .clk_3_N_out(clk_3_wires[53]),
    .clk_3_S_in(clk_3_wires[52]),
    .prog_clk_3_N_out(prog_clk_3_wires[53]),
    .prog_clk_3_S_in(prog_clk_3_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[83]),
    .prog_clk_0_W_in(prog_clk_0_wires[82]),
    .config_enable_S_in(config_enableWires[314]),
    .reset_E_in(resetWires[160]),
    .reset_W_out(resetWires[157]),
    .Test_en_E_in(Test_enWires[160]),
    .Test_en_W_out(Test_enWires[157]),
    .pReset_S_in(pResetWires[314]),
    .chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_25_ccff_tail),
    .chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__15_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__15_ccff_tail)
  );


  cby_1__1_
  cby_2__8_
  (
    .clk_3_N_out(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[56]),
    .prog_clk_3_N_out(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[56]),
    .prog_clk_0_S_out(prog_clk_0_wires[86]),
    .prog_clk_0_W_in(prog_clk_0_wires[85]),
    .config_enable_S_in(config_enableWires[363]),
    .reset_E_in(resetWires[182]),
    .reset_W_out(resetWires[179]),
    .Test_en_E_in(Test_enWires[182]),
    .Test_en_W_out(Test_enWires[179]),
    .pReset_S_in(pResetWires[363]),
    .chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_26_ccff_tail),
    .chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__16_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__16_ccff_tail)
  );


  cby_1__1_
  cby_2__9_
  (
    .clk_3_N_out(clk_3_wires[63]),
    .clk_3_S_in(clk_3_wires[62]),
    .prog_clk_3_N_out(prog_clk_3_wires[63]),
    .prog_clk_3_S_in(prog_clk_3_wires[62]),
    .prog_clk_0_S_out(prog_clk_0_wires[89]),
    .prog_clk_0_W_in(prog_clk_0_wires[88]),
    .config_enable_S_in(config_enableWires[412]),
    .reset_E_in(resetWires[204]),
    .reset_W_out(resetWires[201]),
    .Test_en_E_in(Test_enWires[204]),
    .Test_en_W_out(Test_enWires[201]),
    .pReset_S_in(pResetWires[412]),
    .chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_27_ccff_tail),
    .chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__17_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__17_ccff_tail)
  );


  cby_1__1_
  cby_2__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[95]),
    .prog_clk_0_W_in(prog_clk_0_wires[94]),
    .config_enable_S_in(config_enableWires[510]),
    .reset_E_in(resetWires[248]),
    .reset_W_out(resetWires[245]),
    .Test_en_E_in(Test_enWires[248]),
    .Test_en_W_out(Test_enWires[245]),
    .pReset_S_in(pResetWires[510]),
    .chany_bottom_in(sb_2__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_28_ccff_tail),
    .chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__18_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__18_ccff_tail)
  );


  cby_1__1_
  cby_2__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[100]),
    .prog_clk_0_S_out(prog_clk_0_wires[98]),
    .prog_clk_0_W_in(prog_clk_0_wires[97]),
    .config_enable_S_in(config_enableWires[559]),
    .reset_E_in(resetWires[270]),
    .reset_W_out(resetWires[267]),
    .Test_en_E_in(Test_enWires[270]),
    .Test_en_W_out(Test_enWires[267]),
    .pReset_S_in(pResetWires[559]),
    .chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__1_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__1_ccff_tail),
    .chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__19_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__19_ccff_tail)
  );


  cby_1__1_
  cby_3__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[103]),
    .prog_clk_0_W_in(prog_clk_0_wires[102]),
    .config_enable_S_in(config_enableWires[33]),
    .reset_E_in(resetWires[30]),
    .reset_W_out(resetWires[27]),
    .Test_en_E_in(Test_enWires[30]),
    .Test_en_W_out(Test_enWires[27]),
    .pReset_S_in(pResetWires[33]),
    .chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_30_ccff_tail),
    .chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__20_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__20_ccff_tail)
  );


  cby_1__1_
  cby_3__2_
  (
    .clk_2_S_out(clk_2_wires[30]),
    .clk_2_N_in(clk_2_wires[29]),
    .prog_clk_2_S_out(prog_clk_2_wires[30]),
    .prog_clk_2_N_in(prog_clk_2_wires[29]),
    .prog_clk_0_S_out(prog_clk_0_wires[106]),
    .prog_clk_0_W_in(prog_clk_0_wires[105]),
    .config_enable_S_in(config_enableWires[73]),
    .reset_E_in(resetWires[52]),
    .reset_W_out(resetWires[49]),
    .Test_en_E_in(Test_enWires[52]),
    .Test_en_W_out(Test_enWires[49]),
    .pReset_S_in(pResetWires[73]),
    .chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_31_ccff_tail),
    .chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__21_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__21_ccff_tail)
  );


  cby_1__1_
  cby_3__4_
  (
    .clk_2_S_out(clk_2_wires[41]),
    .clk_2_N_in(clk_2_wires[40]),
    .prog_clk_2_S_out(prog_clk_2_wires[41]),
    .prog_clk_2_N_in(prog_clk_2_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[112]),
    .prog_clk_0_W_in(prog_clk_0_wires[111]),
    .config_enable_S_in(config_enableWires[171]),
    .reset_E_in(resetWires[96]),
    .reset_W_out(resetWires[93]),
    .Test_en_E_in(Test_enWires[96]),
    .Test_en_W_out(Test_enWires[93]),
    .pReset_S_in(pResetWires[171]),
    .chany_bottom_in(sb_1__3__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_32_ccff_tail),
    .chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__22_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__22_ccff_tail)
  );


  cby_1__1_
  cby_3__5_
  (
    .clk_2_N_out(clk_2_wires[39]),
    .clk_2_S_in(clk_2_wires[38]),
    .prog_clk_2_N_out(prog_clk_2_wires[39]),
    .prog_clk_2_S_in(prog_clk_2_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[115]),
    .prog_clk_0_W_in(prog_clk_0_wires[114]),
    .config_enable_S_in(config_enableWires[220]),
    .reset_E_in(resetWires[118]),
    .reset_W_out(resetWires[115]),
    .Test_en_E_in(Test_enWires[118]),
    .Test_en_W_out(Test_enWires[115]),
    .pReset_S_in(pResetWires[220]),
    .chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_33_ccff_tail),
    .chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__23_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__23_ccff_tail)
  );


  cby_1__1_
  cby_3__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[118]),
    .prog_clk_0_W_in(prog_clk_0_wires[117]),
    .config_enable_S_in(config_enableWires[269]),
    .reset_E_in(resetWires[140]),
    .reset_W_out(resetWires[137]),
    .Test_en_E_in(Test_enWires[140]),
    .Test_en_W_out(Test_enWires[137]),
    .pReset_S_in(pResetWires[269]),
    .chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_34_ccff_tail),
    .chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__24_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__24_ccff_tail)
  );


  cby_1__1_
  cby_3__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[121]),
    .prog_clk_0_W_in(prog_clk_0_wires[120]),
    .config_enable_S_in(config_enableWires[318]),
    .reset_E_in(resetWires[162]),
    .reset_W_out(resetWires[159]),
    .Test_en_E_in(Test_enWires[162]),
    .Test_en_W_out(Test_enWires[159]),
    .pReset_S_in(pResetWires[318]),
    .chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_35_ccff_tail),
    .chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__25_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__25_ccff_tail)
  );


  cby_1__1_
  cby_3__8_
  (
    .clk_2_S_out(clk_2_wires[54]),
    .clk_2_N_in(clk_2_wires[53]),
    .prog_clk_2_S_out(prog_clk_2_wires[54]),
    .prog_clk_2_N_in(prog_clk_2_wires[53]),
    .prog_clk_0_S_out(prog_clk_0_wires[124]),
    .prog_clk_0_W_in(prog_clk_0_wires[123]),
    .config_enable_S_in(config_enableWires[367]),
    .reset_E_in(resetWires[184]),
    .reset_W_out(resetWires[181]),
    .Test_en_E_in(Test_enWires[184]),
    .Test_en_W_out(Test_enWires[181]),
    .pReset_S_in(pResetWires[367]),
    .chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_36_ccff_tail),
    .chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__26_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__26_ccff_tail)
  );


  cby_1__1_
  cby_3__9_
  (
    .clk_2_N_out(clk_2_wires[52]),
    .clk_2_S_in(clk_2_wires[51]),
    .prog_clk_2_N_out(prog_clk_2_wires[52]),
    .prog_clk_2_S_in(prog_clk_2_wires[51]),
    .prog_clk_0_S_out(prog_clk_0_wires[127]),
    .prog_clk_0_W_in(prog_clk_0_wires[126]),
    .config_enable_S_in(config_enableWires[416]),
    .reset_E_in(resetWires[206]),
    .reset_W_out(resetWires[203]),
    .Test_en_E_in(Test_enWires[206]),
    .Test_en_W_out(Test_enWires[203]),
    .pReset_S_in(pResetWires[416]),
    .chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_37_ccff_tail),
    .chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__27_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__27_ccff_tail)
  );


  cby_1__1_
  cby_3__11_
  (
    .clk_2_N_out(clk_2_wires[65]),
    .clk_2_S_in(clk_2_wires[64]),
    .prog_clk_2_N_out(prog_clk_2_wires[65]),
    .prog_clk_2_S_in(prog_clk_2_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[133]),
    .prog_clk_0_W_in(prog_clk_0_wires[132]),
    .config_enable_S_in(config_enableWires[514]),
    .reset_E_in(resetWires[250]),
    .reset_W_out(resetWires[247]),
    .Test_en_E_in(Test_enWires[250]),
    .Test_en_W_out(Test_enWires[247]),
    .pReset_S_in(pResetWires[514]),
    .chany_bottom_in(sb_1__3__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_38_ccff_tail),
    .chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__28_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__28_ccff_tail)
  );


  cby_1__1_
  cby_3__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[138]),
    .prog_clk_0_S_out(prog_clk_0_wires[136]),
    .prog_clk_0_W_in(prog_clk_0_wires[135]),
    .config_enable_S_in(config_enableWires[563]),
    .reset_E_in(resetWires[272]),
    .reset_W_out(resetWires[269]),
    .Test_en_E_in(Test_enWires[272]),
    .Test_en_W_out(Test_enWires[269]),
    .pReset_S_in(pResetWires[563]),
    .chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__2_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__2_ccff_tail),
    .chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__29_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__29_ccff_tail)
  );


  cby_1__1_
  cby_4__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[141]),
    .prog_clk_0_W_in(prog_clk_0_wires[140]),
    .config_enable_S_in(config_enableWires[36]),
    .reset_E_in(resetWires[32]),
    .reset_W_out(resetWires[29]),
    .Test_en_E_in(Test_enWires[32]),
    .Test_en_W_out(Test_enWires[29]),
    .pReset_S_in(pResetWires[36]),
    .chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_40_ccff_tail),
    .chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__30_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__30_ccff_tail)
  );


  cby_1__1_
  cby_4__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[144]),
    .prog_clk_0_W_in(prog_clk_0_wires[143]),
    .config_enable_S_in(config_enableWires[77]),
    .reset_E_in(resetWires[54]),
    .reset_W_out(resetWires[51]),
    .Test_en_E_in(Test_enWires[54]),
    .Test_en_W_out(Test_enWires[51]),
    .pReset_S_in(pResetWires[77]),
    .chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_41_ccff_tail),
    .chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__31_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__31_ccff_tail)
  );


  cby_1__1_
  cby_4__4_
  (
    .clk_3_S_out(clk_3_wires[21]),
    .clk_3_N_in(clk_3_wires[20]),
    .prog_clk_3_S_out(prog_clk_3_wires[21]),
    .prog_clk_3_N_in(prog_clk_3_wires[20]),
    .prog_clk_0_S_out(prog_clk_0_wires[150]),
    .prog_clk_0_W_in(prog_clk_0_wires[149]),
    .config_enable_S_in(config_enableWires[175]),
    .reset_E_in(resetWires[98]),
    .reset_W_out(resetWires[95]),
    .Test_en_E_in(Test_enWires[98]),
    .Test_en_W_out(Test_enWires[95]),
    .pReset_S_in(pResetWires[175]),
    .chany_bottom_in(sb_2__3__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_42_ccff_tail),
    .chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__32_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__32_ccff_tail)
  );


  cby_1__1_
  cby_4__5_
  (
    .clk_3_S_out(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[14]),
    .prog_clk_3_S_out(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[14]),
    .prog_clk_0_S_out(prog_clk_0_wires[153]),
    .prog_clk_0_W_in(prog_clk_0_wires[152]),
    .config_enable_S_in(config_enableWires[224]),
    .reset_E_in(resetWires[120]),
    .reset_W_out(resetWires[117]),
    .Test_en_E_in(Test_enWires[120]),
    .Test_en_W_out(Test_enWires[117]),
    .pReset_S_in(pResetWires[224]),
    .chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_43_ccff_tail),
    .chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__33_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__33_ccff_tail)
  );


  cby_1__1_
  cby_4__6_
  (
    .clk_3_S_out(clk_3_wires[11]),
    .clk_3_N_in(clk_3_wires[10]),
    .prog_clk_3_S_out(prog_clk_3_wires[11]),
    .prog_clk_3_N_in(prog_clk_3_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[156]),
    .prog_clk_0_W_in(prog_clk_0_wires[155]),
    .config_enable_S_in(config_enableWires[273]),
    .reset_E_in(resetWires[142]),
    .reset_W_out(resetWires[139]),
    .Test_en_E_in(Test_enWires[142]),
    .Test_en_W_out(Test_enWires[139]),
    .pReset_S_in(pResetWires[273]),
    .chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_44_ccff_tail),
    .chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__34_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__34_ccff_tail)
  );


  cby_1__1_
  cby_4__7_
  (
    .clk_3_N_out(clk_3_wires[9]),
    .clk_3_S_in(clk_3_wires[8]),
    .prog_clk_3_N_out(prog_clk_3_wires[9]),
    .prog_clk_3_S_in(prog_clk_3_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[159]),
    .prog_clk_0_W_in(prog_clk_0_wires[158]),
    .config_enable_S_in(config_enableWires[322]),
    .reset_E_in(resetWires[164]),
    .reset_W_out(resetWires[161]),
    .Test_en_E_in(Test_enWires[164]),
    .Test_en_W_out(Test_enWires[161]),
    .pReset_S_in(pResetWires[322]),
    .chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_45_ccff_tail),
    .chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__35_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__35_ccff_tail)
  );


  cby_1__1_
  cby_4__8_
  (
    .clk_3_N_out(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[12]),
    .prog_clk_3_N_out(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[162]),
    .prog_clk_0_W_in(prog_clk_0_wires[161]),
    .config_enable_S_in(config_enableWires[371]),
    .reset_E_in(resetWires[186]),
    .reset_W_out(resetWires[183]),
    .Test_en_E_in(Test_enWires[186]),
    .Test_en_W_out(Test_enWires[183]),
    .pReset_S_in(pResetWires[371]),
    .chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_46_ccff_tail),
    .chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__36_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__36_ccff_tail)
  );


  cby_1__1_
  cby_4__9_
  (
    .clk_3_N_out(clk_3_wires[19]),
    .clk_3_S_in(clk_3_wires[18]),
    .prog_clk_3_N_out(prog_clk_3_wires[19]),
    .prog_clk_3_S_in(prog_clk_3_wires[18]),
    .prog_clk_0_S_out(prog_clk_0_wires[165]),
    .prog_clk_0_W_in(prog_clk_0_wires[164]),
    .config_enable_S_in(config_enableWires[420]),
    .reset_E_in(resetWires[208]),
    .reset_W_out(resetWires[205]),
    .Test_en_E_in(Test_enWires[208]),
    .Test_en_W_out(Test_enWires[205]),
    .pReset_S_in(pResetWires[420]),
    .chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_47_ccff_tail),
    .chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__37_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__37_ccff_tail)
  );


  cby_1__1_
  cby_4__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[171]),
    .prog_clk_0_W_in(prog_clk_0_wires[170]),
    .config_enable_S_in(config_enableWires[518]),
    .reset_E_in(resetWires[252]),
    .reset_W_out(resetWires[249]),
    .Test_en_E_in(Test_enWires[252]),
    .Test_en_W_out(Test_enWires[249]),
    .pReset_S_in(pResetWires[518]),
    .chany_bottom_in(sb_2__3__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_48_ccff_tail),
    .chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__38_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__38_ccff_tail)
  );


  cby_1__1_
  cby_4__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[176]),
    .prog_clk_0_S_out(prog_clk_0_wires[174]),
    .prog_clk_0_W_in(prog_clk_0_wires[173]),
    .config_enable_S_in(config_enableWires[567]),
    .reset_E_in(resetWires[274]),
    .reset_W_out(resetWires[271]),
    .Test_en_E_in(Test_enWires[274]),
    .Test_en_W_out(Test_enWires[271]),
    .pReset_S_in(pResetWires[567]),
    .chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__3_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__3_ccff_tail),
    .chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__39_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__39_ccff_tail)
  );


  cby_1__1_
  cby_5__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[179]),
    .prog_clk_0_W_in(prog_clk_0_wires[178]),
    .config_enable_S_in(config_enableWires[39]),
    .reset_E_in(resetWires[34]),
    .reset_W_out(resetWires[31]),
    .Test_en_E_in(Test_enWires[34]),
    .Test_en_W_out(Test_enWires[31]),
    .pReset_S_in(pResetWires[39]),
    .chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_50_ccff_tail),
    .chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__40_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__40_ccff_tail)
  );


  cby_1__1_
  cby_5__2_
  (
    .clk_2_S_out(clk_2_wires[32]),
    .clk_2_N_in(clk_2_wires[31]),
    .prog_clk_2_S_out(prog_clk_2_wires[32]),
    .prog_clk_2_N_in(prog_clk_2_wires[31]),
    .prog_clk_0_S_out(prog_clk_0_wires[182]),
    .prog_clk_0_W_in(prog_clk_0_wires[181]),
    .config_enable_S_in(config_enableWires[81]),
    .reset_E_in(resetWires[56]),
    .reset_W_out(resetWires[53]),
    .Test_en_E_in(Test_enWires[56]),
    .Test_en_W_out(Test_enWires[53]),
    .pReset_S_in(pResetWires[81]),
    .chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_51_ccff_tail),
    .chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__41_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__41_ccff_tail)
  );


  cby_1__1_
  cby_5__4_
  (
    .clk_2_S_out(clk_2_wires[45]),
    .clk_2_N_in(clk_2_wires[44]),
    .prog_clk_2_S_out(prog_clk_2_wires[45]),
    .prog_clk_2_N_in(prog_clk_2_wires[44]),
    .prog_clk_0_S_out(prog_clk_0_wires[188]),
    .prog_clk_0_W_in(prog_clk_0_wires[187]),
    .config_enable_S_in(config_enableWires[179]),
    .reset_E_in(resetWires[100]),
    .reset_W_out(resetWires[97]),
    .Test_en_E_in(Test_enWires[100]),
    .Test_en_W_out(Test_enWires[97]),
    .pReset_S_in(pResetWires[179]),
    .chany_bottom_in(sb_1__3__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_52_ccff_tail),
    .chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__42_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__42_ccff_tail)
  );


  cby_1__1_
  cby_5__5_
  (
    .clk_2_N_out(clk_2_wires[43]),
    .clk_2_S_in(clk_2_wires[42]),
    .prog_clk_2_N_out(prog_clk_2_wires[43]),
    .prog_clk_2_S_in(prog_clk_2_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[191]),
    .prog_clk_0_W_in(prog_clk_0_wires[190]),
    .config_enable_S_in(config_enableWires[228]),
    .reset_E_in(resetWires[122]),
    .reset_W_out(resetWires[119]),
    .Test_en_E_in(Test_enWires[122]),
    .Test_en_W_out(Test_enWires[119]),
    .pReset_S_in(pResetWires[228]),
    .chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_53_ccff_tail),
    .chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__43_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__43_ccff_tail)
  );


  cby_1__1_
  cby_5__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[194]),
    .prog_clk_0_W_in(prog_clk_0_wires[193]),
    .config_enable_S_in(config_enableWires[277]),
    .reset_E_in(resetWires[144]),
    .reset_W_out(resetWires[141]),
    .Test_en_E_in(Test_enWires[144]),
    .Test_en_W_out(Test_enWires[141]),
    .pReset_S_in(pResetWires[277]),
    .chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_54_ccff_tail),
    .chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__44_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__44_ccff_tail)
  );


  cby_1__1_
  cby_5__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[197]),
    .prog_clk_0_W_in(prog_clk_0_wires[196]),
    .config_enable_S_in(config_enableWires[326]),
    .reset_E_in(resetWires[166]),
    .reset_W_out(resetWires[163]),
    .Test_en_E_in(Test_enWires[166]),
    .Test_en_W_out(Test_enWires[163]),
    .pReset_S_in(pResetWires[326]),
    .chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_55_ccff_tail),
    .chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__45_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__45_ccff_tail)
  );


  cby_1__1_
  cby_5__8_
  (
    .clk_2_S_out(clk_2_wires[58]),
    .clk_2_N_in(clk_2_wires[57]),
    .prog_clk_2_S_out(prog_clk_2_wires[58]),
    .prog_clk_2_N_in(prog_clk_2_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[200]),
    .prog_clk_0_W_in(prog_clk_0_wires[199]),
    .config_enable_S_in(config_enableWires[375]),
    .reset_E_in(resetWires[188]),
    .reset_W_out(resetWires[185]),
    .Test_en_E_in(Test_enWires[188]),
    .Test_en_W_out(Test_enWires[185]),
    .pReset_S_in(pResetWires[375]),
    .chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_56_ccff_tail),
    .chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__46_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__46_ccff_tail)
  );


  cby_1__1_
  cby_5__9_
  (
    .clk_2_N_out(clk_2_wires[56]),
    .clk_2_S_in(clk_2_wires[55]),
    .prog_clk_2_N_out(prog_clk_2_wires[56]),
    .prog_clk_2_S_in(prog_clk_2_wires[55]),
    .prog_clk_0_S_out(prog_clk_0_wires[203]),
    .prog_clk_0_W_in(prog_clk_0_wires[202]),
    .config_enable_S_in(config_enableWires[424]),
    .reset_E_in(resetWires[210]),
    .reset_W_out(resetWires[207]),
    .Test_en_E_in(Test_enWires[210]),
    .Test_en_W_out(Test_enWires[207]),
    .pReset_S_in(pResetWires[424]),
    .chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_57_ccff_tail),
    .chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__47_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__47_ccff_tail)
  );


  cby_1__1_
  cby_5__11_
  (
    .clk_2_N_out(clk_2_wires[67]),
    .clk_2_S_in(clk_2_wires[66]),
    .prog_clk_2_N_out(prog_clk_2_wires[67]),
    .prog_clk_2_S_in(prog_clk_2_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[209]),
    .prog_clk_0_W_in(prog_clk_0_wires[208]),
    .config_enable_S_in(config_enableWires[522]),
    .reset_E_in(resetWires[254]),
    .reset_W_out(resetWires[251]),
    .Test_en_E_in(Test_enWires[254]),
    .Test_en_W_out(Test_enWires[251]),
    .pReset_S_in(pResetWires[522]),
    .chany_bottom_in(sb_1__3__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_58_ccff_tail),
    .chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__48_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__48_ccff_tail)
  );


  cby_1__1_
  cby_5__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[214]),
    .prog_clk_0_S_out(prog_clk_0_wires[212]),
    .prog_clk_0_W_in(prog_clk_0_wires[211]),
    .config_enable_S_in(config_enableWires[571]),
    .reset_E_in(resetWires[276]),
    .reset_W_out(resetWires[273]),
    .Test_en_E_in(Test_enWires[276]),
    .Test_en_W_out(Test_enWires[273]),
    .pReset_S_in(pResetWires[571]),
    .chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__4_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__4_ccff_tail),
    .chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__49_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__49_ccff_tail)
  );


  cby_1__1_
  cby_6__1_
  (
    .clk_3_S_in(clk_3_wires[90]),
    .clk_3_N_out(clk_3_wires[89]),
    .prog_clk_3_S_in(prog_clk_3_wires[90]),
    .prog_clk_3_N_out(prog_clk_3_wires[89]),
    .prog_clk_0_S_out(prog_clk_0_wires[217]),
    .prog_clk_0_W_in(prog_clk_0_wires[216]),
    .config_enable_N_out(config_enableWires[2]),
    .config_enable_S_in(config_enableWires[42]),
    .reset_E_out(resetWires[35]),
    .reset_W_out(resetWires[33]),
    .reset_N_out(resetWires[2]),
    .reset_S_in(resetWires[1]),
    .Test_en_E_out(Test_enWires[35]),
    .Test_en_W_out(Test_enWires[33]),
    .Test_en_N_out(Test_enWires[2]),
    .Test_en_S_in(Test_enWires[1]),
    .pReset_N_out(pResetWires[2]),
    .pReset_S_in(pResetWires[42]),
    .chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_60_ccff_tail),
    .chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__50_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__50_ccff_tail)
  );


  cby_1__1_
  cby_6__2_
  (
    .clk_3_S_in(clk_3_wires[92]),
    .clk_3_N_out(clk_3_wires[91]),
    .prog_clk_3_S_in(prog_clk_3_wires[92]),
    .prog_clk_3_N_out(prog_clk_3_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[220]),
    .prog_clk_0_W_in(prog_clk_0_wires[219]),
    .config_enable_N_out(config_enableWires[4]),
    .config_enable_S_in(config_enableWires[85]),
    .reset_E_out(resetWires[57]),
    .reset_W_out(resetWires[55]),
    .reset_N_out(resetWires[4]),
    .reset_S_in(resetWires[3]),
    .Test_en_E_out(Test_enWires[57]),
    .Test_en_W_out(Test_enWires[55]),
    .Test_en_N_out(Test_enWires[4]),
    .Test_en_S_in(Test_enWires[3]),
    .pReset_N_out(pResetWires[4]),
    .pReset_S_in(pResetWires[85]),
    .chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_61_ccff_tail),
    .chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__51_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__51_ccff_tail)
  );


  cby_1__1_
  cby_6__4_
  (
    .clk_3_S_in(clk_3_wires[96]),
    .clk_3_N_out(clk_3_wires[95]),
    .prog_clk_3_S_in(prog_clk_3_wires[96]),
    .prog_clk_3_N_out(prog_clk_3_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[226]),
    .prog_clk_0_W_in(prog_clk_0_wires[225]),
    .config_enable_N_out(config_enableWires[8]),
    .config_enable_S_in(config_enableWires[183]),
    .reset_E_out(resetWires[101]),
    .reset_W_out(resetWires[99]),
    .reset_N_out(resetWires[8]),
    .reset_S_in(resetWires[7]),
    .Test_en_E_out(Test_enWires[101]),
    .Test_en_W_out(Test_enWires[99]),
    .Test_en_N_out(Test_enWires[8]),
    .Test_en_S_in(Test_enWires[7]),
    .pReset_N_out(pResetWires[8]),
    .pReset_S_in(pResetWires[183]),
    .chany_bottom_in(sb_2__3__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_62_ccff_tail),
    .chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__52_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__52_ccff_tail)
  );


  cby_1__1_
  cby_6__5_
  (
    .clk_3_S_in(clk_3_wires[98]),
    .clk_3_N_out(clk_3_wires[97]),
    .prog_clk_3_S_in(prog_clk_3_wires[98]),
    .prog_clk_3_N_out(prog_clk_3_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[229]),
    .prog_clk_0_W_in(prog_clk_0_wires[228]),
    .config_enable_N_out(config_enableWires[10]),
    .config_enable_S_in(config_enableWires[232]),
    .reset_E_out(resetWires[123]),
    .reset_W_out(resetWires[121]),
    .reset_N_out(resetWires[10]),
    .reset_S_in(resetWires[9]),
    .Test_en_E_out(Test_enWires[123]),
    .Test_en_W_out(Test_enWires[121]),
    .Test_en_N_out(Test_enWires[10]),
    .Test_en_S_in(Test_enWires[9]),
    .pReset_N_out(pResetWires[10]),
    .pReset_S_in(pResetWires[232]),
    .chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_63_ccff_tail),
    .chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__53_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__53_ccff_tail)
  );


  cby_1__1_
  cby_6__6_
  (
    .clk_3_S_in(clk_3_wires[100]),
    .clk_3_N_out(clk_3_wires[99]),
    .prog_clk_3_S_in(prog_clk_3_wires[100]),
    .prog_clk_3_N_out(prog_clk_3_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[232]),
    .prog_clk_0_W_in(prog_clk_0_wires[231]),
    .config_enable_N_out(config_enableWires[12]),
    .config_enable_S_in(config_enableWires[281]),
    .reset_E_out(resetWires[145]),
    .reset_W_out(resetWires[143]),
    .reset_N_out(resetWires[12]),
    .reset_S_in(resetWires[11]),
    .Test_en_E_out(Test_enWires[145]),
    .Test_en_W_out(Test_enWires[143]),
    .Test_en_N_out(Test_enWires[12]),
    .Test_en_S_in(Test_enWires[11]),
    .pReset_N_out(pResetWires[12]),
    .pReset_S_in(pResetWires[281]),
    .chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_64_ccff_tail),
    .chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__54_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__54_ccff_tail)
  );


  cby_1__1_
  cby_6__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[235]),
    .prog_clk_0_W_in(prog_clk_0_wires[234]),
    .config_enable_N_out(config_enableWires[14]),
    .config_enable_S_in(config_enableWires[330]),
    .reset_E_out(resetWires[167]),
    .reset_W_out(resetWires[165]),
    .reset_N_out(resetWires[14]),
    .reset_S_in(resetWires[13]),
    .Test_en_E_out(Test_enWires[167]),
    .Test_en_W_out(Test_enWires[165]),
    .Test_en_N_out(Test_enWires[14]),
    .Test_en_S_in(Test_enWires[13]),
    .pReset_N_out(pResetWires[14]),
    .pReset_S_in(pResetWires[330]),
    .chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_65_ccff_tail),
    .chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__55_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__55_ccff_tail)
  );


  cby_1__1_
  cby_6__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[238]),
    .prog_clk_0_W_in(prog_clk_0_wires[237]),
    .config_enable_N_out(config_enableWires[16]),
    .config_enable_S_in(config_enableWires[379]),
    .reset_E_out(resetWires[189]),
    .reset_W_out(resetWires[187]),
    .reset_N_out(resetWires[16]),
    .reset_S_in(resetWires[15]),
    .Test_en_E_out(Test_enWires[189]),
    .Test_en_W_out(Test_enWires[187]),
    .Test_en_N_out(Test_enWires[16]),
    .Test_en_S_in(Test_enWires[15]),
    .pReset_N_out(pResetWires[16]),
    .pReset_S_in(pResetWires[379]),
    .chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_66_ccff_tail),
    .chany_bottom_out(cby_1__1__56_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__56_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__56_ccff_tail)
  );


  cby_1__1_
  cby_6__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[241]),
    .prog_clk_0_W_in(prog_clk_0_wires[240]),
    .config_enable_N_out(config_enableWires[18]),
    .config_enable_S_in(config_enableWires[428]),
    .reset_E_out(resetWires[211]),
    .reset_W_out(resetWires[209]),
    .reset_N_out(resetWires[18]),
    .reset_S_in(resetWires[17]),
    .Test_en_E_out(Test_enWires[211]),
    .Test_en_W_out(Test_enWires[209]),
    .Test_en_N_out(Test_enWires[18]),
    .Test_en_S_in(Test_enWires[17]),
    .pReset_N_out(pResetWires[18]),
    .pReset_S_in(pResetWires[428]),
    .chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_67_ccff_tail),
    .chany_bottom_out(cby_1__1__57_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__57_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__57_ccff_tail)
  );


  cby_1__1_
  cby_6__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[247]),
    .prog_clk_0_W_in(prog_clk_0_wires[246]),
    .config_enable_N_out(config_enableWires[22]),
    .config_enable_S_in(config_enableWires[526]),
    .reset_E_out(resetWires[255]),
    .reset_W_out(resetWires[253]),
    .reset_N_out(resetWires[22]),
    .reset_S_in(resetWires[21]),
    .Test_en_E_out(Test_enWires[255]),
    .Test_en_W_out(Test_enWires[253]),
    .Test_en_N_out(Test_enWires[22]),
    .Test_en_S_in(Test_enWires[21]),
    .pReset_N_out(pResetWires[22]),
    .pReset_S_in(pResetWires[526]),
    .chany_bottom_in(sb_2__3__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_68_ccff_tail),
    .chany_bottom_out(cby_1__1__58_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__58_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__58_ccff_tail)
  );


  cby_1__1_
  cby_6__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[252]),
    .prog_clk_0_S_out(prog_clk_0_wires[250]),
    .prog_clk_0_W_in(prog_clk_0_wires[249]),
    .config_enable_N_out(config_enableWires[24]),
    .config_enable_S_in(config_enableWires[575]),
    .reset_E_out(resetWires[277]),
    .reset_W_out(resetWires[275]),
    .reset_S_in(resetWires[23]),
    .Test_en_E_out(Test_enWires[277]),
    .Test_en_W_out(Test_enWires[275]),
    .Test_en_S_in(Test_enWires[23]),
    .pReset_N_out(pResetWires[24]),
    .pReset_S_in(pResetWires[575]),
    .chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__5_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__5_ccff_tail),
    .chany_bottom_out(cby_1__1__59_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__59_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__59_ccff_tail)
  );


  cby_1__1_
  cby_7__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[255]),
    .prog_clk_0_W_in(prog_clk_0_wires[254]),
    .config_enable_S_in(config_enableWires[45]),
    .reset_E_out(resetWires[37]),
    .reset_W_in(resetWires[36]),
    .Test_en_E_out(Test_enWires[37]),
    .Test_en_W_in(Test_enWires[36]),
    .pReset_S_in(pResetWires[45]),
    .chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_70_ccff_tail),
    .chany_bottom_out(cby_1__1__60_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__60_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__60_ccff_tail)
  );


  cby_1__1_
  cby_7__2_
  (
    .clk_2_S_out(clk_2_wires[74]),
    .clk_2_N_in(clk_2_wires[73]),
    .prog_clk_2_S_out(prog_clk_2_wires[74]),
    .prog_clk_2_N_in(prog_clk_2_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[258]),
    .prog_clk_0_W_in(prog_clk_0_wires[257]),
    .config_enable_S_in(config_enableWires[89]),
    .reset_E_out(resetWires[59]),
    .reset_W_in(resetWires[58]),
    .Test_en_E_out(Test_enWires[59]),
    .Test_en_W_in(Test_enWires[58]),
    .pReset_S_in(pResetWires[89]),
    .chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_71_ccff_tail),
    .chany_bottom_out(cby_1__1__61_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__61_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__61_ccff_tail)
  );


  cby_1__1_
  cby_7__4_
  (
    .clk_2_S_out(clk_2_wires[85]),
    .clk_2_N_in(clk_2_wires[84]),
    .prog_clk_2_S_out(prog_clk_2_wires[85]),
    .prog_clk_2_N_in(prog_clk_2_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[264]),
    .prog_clk_0_W_in(prog_clk_0_wires[263]),
    .config_enable_S_in(config_enableWires[187]),
    .reset_E_out(resetWires[103]),
    .reset_W_in(resetWires[102]),
    .Test_en_E_out(Test_enWires[103]),
    .Test_en_W_in(Test_enWires[102]),
    .pReset_S_in(pResetWires[187]),
    .chany_bottom_in(sb_1__3__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_72_ccff_tail),
    .chany_bottom_out(cby_1__1__62_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__62_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__62_ccff_tail)
  );


  cby_1__1_
  cby_7__5_
  (
    .clk_2_N_out(clk_2_wires[83]),
    .clk_2_S_in(clk_2_wires[82]),
    .prog_clk_2_N_out(prog_clk_2_wires[83]),
    .prog_clk_2_S_in(prog_clk_2_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[267]),
    .prog_clk_0_W_in(prog_clk_0_wires[266]),
    .config_enable_S_in(config_enableWires[236]),
    .reset_E_out(resetWires[125]),
    .reset_W_in(resetWires[124]),
    .Test_en_E_out(Test_enWires[125]),
    .Test_en_W_in(Test_enWires[124]),
    .pReset_S_in(pResetWires[236]),
    .chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_73_ccff_tail),
    .chany_bottom_out(cby_1__1__63_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__63_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__63_ccff_tail)
  );


  cby_1__1_
  cby_7__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[270]),
    .prog_clk_0_W_in(prog_clk_0_wires[269]),
    .config_enable_S_in(config_enableWires[285]),
    .reset_E_out(resetWires[147]),
    .reset_W_in(resetWires[146]),
    .Test_en_E_out(Test_enWires[147]),
    .Test_en_W_in(Test_enWires[146]),
    .pReset_S_in(pResetWires[285]),
    .chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_74_ccff_tail),
    .chany_bottom_out(cby_1__1__64_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__64_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__64_ccff_tail)
  );


  cby_1__1_
  cby_7__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[273]),
    .prog_clk_0_W_in(prog_clk_0_wires[272]),
    .config_enable_S_in(config_enableWires[334]),
    .reset_E_out(resetWires[169]),
    .reset_W_in(resetWires[168]),
    .Test_en_E_out(Test_enWires[169]),
    .Test_en_W_in(Test_enWires[168]),
    .pReset_S_in(pResetWires[334]),
    .chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_75_ccff_tail),
    .chany_bottom_out(cby_1__1__65_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__65_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__65_ccff_tail)
  );


  cby_1__1_
  cby_7__8_
  (
    .clk_2_S_out(clk_2_wires[98]),
    .clk_2_N_in(clk_2_wires[97]),
    .prog_clk_2_S_out(prog_clk_2_wires[98]),
    .prog_clk_2_N_in(prog_clk_2_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[276]),
    .prog_clk_0_W_in(prog_clk_0_wires[275]),
    .config_enable_S_in(config_enableWires[383]),
    .reset_E_out(resetWires[191]),
    .reset_W_in(resetWires[190]),
    .Test_en_E_out(Test_enWires[191]),
    .Test_en_W_in(Test_enWires[190]),
    .pReset_S_in(pResetWires[383]),
    .chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_76_ccff_tail),
    .chany_bottom_out(cby_1__1__66_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__66_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__66_ccff_tail)
  );


  cby_1__1_
  cby_7__9_
  (
    .clk_2_N_out(clk_2_wires[96]),
    .clk_2_S_in(clk_2_wires[95]),
    .prog_clk_2_N_out(prog_clk_2_wires[96]),
    .prog_clk_2_S_in(prog_clk_2_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[279]),
    .prog_clk_0_W_in(prog_clk_0_wires[278]),
    .config_enable_S_in(config_enableWires[432]),
    .reset_E_out(resetWires[213]),
    .reset_W_in(resetWires[212]),
    .Test_en_E_out(Test_enWires[213]),
    .Test_en_W_in(Test_enWires[212]),
    .pReset_S_in(pResetWires[432]),
    .chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_77_ccff_tail),
    .chany_bottom_out(cby_1__1__67_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__67_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__67_ccff_tail)
  );


  cby_1__1_
  cby_7__11_
  (
    .clk_2_N_out(clk_2_wires[109]),
    .clk_2_S_in(clk_2_wires[108]),
    .prog_clk_2_N_out(prog_clk_2_wires[109]),
    .prog_clk_2_S_in(prog_clk_2_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[285]),
    .prog_clk_0_W_in(prog_clk_0_wires[284]),
    .config_enable_S_in(config_enableWires[530]),
    .reset_E_out(resetWires[257]),
    .reset_W_in(resetWires[256]),
    .Test_en_E_out(Test_enWires[257]),
    .Test_en_W_in(Test_enWires[256]),
    .pReset_S_in(pResetWires[530]),
    .chany_bottom_in(sb_1__3__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_78_ccff_tail),
    .chany_bottom_out(cby_1__1__68_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__68_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__68_ccff_tail)
  );


  cby_1__1_
  cby_7__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[290]),
    .prog_clk_0_S_out(prog_clk_0_wires[288]),
    .prog_clk_0_W_in(prog_clk_0_wires[287]),
    .config_enable_S_in(config_enableWires[579]),
    .reset_E_out(resetWires[279]),
    .reset_W_in(resetWires[278]),
    .Test_en_E_out(Test_enWires[279]),
    .Test_en_W_in(Test_enWires[278]),
    .pReset_S_in(pResetWires[579]),
    .chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__6_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__6_ccff_tail),
    .chany_bottom_out(cby_1__1__69_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__69_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__69_ccff_tail)
  );


  cby_1__1_
  cby_8__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[293]),
    .prog_clk_0_W_in(prog_clk_0_wires[292]),
    .config_enable_S_in(config_enableWires[48]),
    .reset_E_out(resetWires[39]),
    .reset_W_in(resetWires[38]),
    .Test_en_E_out(Test_enWires[39]),
    .Test_en_W_in(Test_enWires[38]),
    .pReset_S_in(pResetWires[48]),
    .chany_bottom_in(sb_1__0__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__49_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_80_ccff_tail),
    .chany_bottom_out(cby_1__1__70_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__70_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__70_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__70_ccff_tail)
  );


  cby_1__1_
  cby_8__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[296]),
    .prog_clk_0_W_in(prog_clk_0_wires[295]),
    .config_enable_S_in(config_enableWires[93]),
    .reset_E_out(resetWires[61]),
    .reset_W_in(resetWires[60]),
    .Test_en_E_out(Test_enWires[61]),
    .Test_en_W_in(Test_enWires[60]),
    .pReset_S_in(pResetWires[93]),
    .chany_bottom_in(sb_1__1__49_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_81_ccff_tail),
    .chany_bottom_out(cby_1__1__71_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__71_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__71_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__71_ccff_tail)
  );


  cby_1__1_
  cby_8__4_
  (
    .clk_3_S_out(clk_3_wires[39]),
    .clk_3_N_in(clk_3_wires[38]),
    .prog_clk_3_S_out(prog_clk_3_wires[39]),
    .prog_clk_3_N_in(prog_clk_3_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[302]),
    .prog_clk_0_W_in(prog_clk_0_wires[301]),
    .config_enable_S_in(config_enableWires[191]),
    .reset_E_out(resetWires[105]),
    .reset_W_in(resetWires[104]),
    .Test_en_E_out(Test_enWires[105]),
    .Test_en_W_in(Test_enWires[104]),
    .pReset_S_in(pResetWires[191]),
    .chany_bottom_in(sb_2__3__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__50_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_82_ccff_tail),
    .chany_bottom_out(cby_1__1__72_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__72_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__72_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__72_ccff_tail)
  );


  cby_1__1_
  cby_8__5_
  (
    .clk_3_S_out(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[32]),
    .prog_clk_3_S_out(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[305]),
    .prog_clk_0_W_in(prog_clk_0_wires[304]),
    .config_enable_S_in(config_enableWires[240]),
    .reset_E_out(resetWires[127]),
    .reset_W_in(resetWires[126]),
    .Test_en_E_out(Test_enWires[127]),
    .Test_en_W_in(Test_enWires[126]),
    .pReset_S_in(pResetWires[240]),
    .chany_bottom_in(sb_1__1__50_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__51_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_83_ccff_tail),
    .chany_bottom_out(cby_1__1__73_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__73_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__73_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__73_ccff_tail)
  );


  cby_1__1_
  cby_8__6_
  (
    .clk_3_S_out(clk_3_wires[29]),
    .clk_3_N_in(clk_3_wires[28]),
    .prog_clk_3_S_out(prog_clk_3_wires[29]),
    .prog_clk_3_N_in(prog_clk_3_wires[28]),
    .prog_clk_0_S_out(prog_clk_0_wires[308]),
    .prog_clk_0_W_in(prog_clk_0_wires[307]),
    .config_enable_S_in(config_enableWires[289]),
    .reset_E_out(resetWires[149]),
    .reset_W_in(resetWires[148]),
    .Test_en_E_out(Test_enWires[149]),
    .Test_en_W_in(Test_enWires[148]),
    .pReset_S_in(pResetWires[289]),
    .chany_bottom_in(sb_1__1__51_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__52_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_84_ccff_tail),
    .chany_bottom_out(cby_1__1__74_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__74_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__74_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__74_ccff_tail)
  );


  cby_1__1_
  cby_8__7_
  (
    .clk_3_N_out(clk_3_wires[27]),
    .clk_3_S_in(clk_3_wires[26]),
    .prog_clk_3_N_out(prog_clk_3_wires[27]),
    .prog_clk_3_S_in(prog_clk_3_wires[26]),
    .prog_clk_0_S_out(prog_clk_0_wires[311]),
    .prog_clk_0_W_in(prog_clk_0_wires[310]),
    .config_enable_S_in(config_enableWires[338]),
    .reset_E_out(resetWires[171]),
    .reset_W_in(resetWires[170]),
    .Test_en_E_out(Test_enWires[171]),
    .Test_en_W_in(Test_enWires[170]),
    .pReset_S_in(pResetWires[338]),
    .chany_bottom_in(sb_1__1__52_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__53_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_85_ccff_tail),
    .chany_bottom_out(cby_1__1__75_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__75_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__75_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__75_ccff_tail)
  );


  cby_1__1_
  cby_8__8_
  (
    .clk_3_N_out(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[30]),
    .prog_clk_3_N_out(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[30]),
    .prog_clk_0_S_out(prog_clk_0_wires[314]),
    .prog_clk_0_W_in(prog_clk_0_wires[313]),
    .config_enable_S_in(config_enableWires[387]),
    .reset_E_out(resetWires[193]),
    .reset_W_in(resetWires[192]),
    .Test_en_E_out(Test_enWires[193]),
    .Test_en_W_in(Test_enWires[192]),
    .pReset_S_in(pResetWires[387]),
    .chany_bottom_in(sb_1__1__53_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__54_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_86_ccff_tail),
    .chany_bottom_out(cby_1__1__76_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__76_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__76_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__76_ccff_tail)
  );


  cby_1__1_
  cby_8__9_
  (
    .clk_3_N_out(clk_3_wires[37]),
    .clk_3_S_in(clk_3_wires[36]),
    .prog_clk_3_N_out(prog_clk_3_wires[37]),
    .prog_clk_3_S_in(prog_clk_3_wires[36]),
    .prog_clk_0_S_out(prog_clk_0_wires[317]),
    .prog_clk_0_W_in(prog_clk_0_wires[316]),
    .config_enable_S_in(config_enableWires[436]),
    .reset_E_out(resetWires[215]),
    .reset_W_in(resetWires[214]),
    .Test_en_E_out(Test_enWires[215]),
    .Test_en_W_in(Test_enWires[214]),
    .pReset_S_in(pResetWires[436]),
    .chany_bottom_in(sb_1__1__54_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_87_ccff_tail),
    .chany_bottom_out(cby_1__1__77_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__77_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__77_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__77_ccff_tail)
  );


  cby_1__1_
  cby_8__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[323]),
    .prog_clk_0_W_in(prog_clk_0_wires[322]),
    .config_enable_S_in(config_enableWires[534]),
    .reset_E_out(resetWires[259]),
    .reset_W_in(resetWires[258]),
    .Test_en_E_out(Test_enWires[259]),
    .Test_en_W_in(Test_enWires[258]),
    .pReset_S_in(pResetWires[534]),
    .chany_bottom_in(sb_2__3__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__55_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_88_ccff_tail),
    .chany_bottom_out(cby_1__1__78_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__78_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__78_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__78_ccff_tail)
  );


  cby_1__1_
  cby_8__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[328]),
    .prog_clk_0_S_out(prog_clk_0_wires[326]),
    .prog_clk_0_W_in(prog_clk_0_wires[325]),
    .config_enable_S_in(config_enableWires[583]),
    .reset_E_out(resetWires[281]),
    .reset_W_in(resetWires[280]),
    .Test_en_E_out(Test_enWires[281]),
    .Test_en_W_in(Test_enWires[280]),
    .pReset_S_in(pResetWires[583]),
    .chany_bottom_in(sb_1__1__55_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__7_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__7_ccff_tail),
    .chany_bottom_out(cby_1__1__79_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__79_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__79_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__79_ccff_tail)
  );


  cby_1__1_
  cby_9__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[331]),
    .prog_clk_0_W_in(prog_clk_0_wires[330]),
    .config_enable_S_in(config_enableWires[51]),
    .reset_E_out(resetWires[41]),
    .reset_W_in(resetWires[40]),
    .Test_en_E_out(Test_enWires[41]),
    .Test_en_W_in(Test_enWires[40]),
    .pReset_S_in(pResetWires[51]),
    .chany_bottom_in(sb_1__0__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__56_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_90_ccff_tail),
    .chany_bottom_out(cby_1__1__80_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__80_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__80_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__80_ccff_tail)
  );


  cby_1__1_
  cby_9__2_
  (
    .clk_2_S_out(clk_2_wires[76]),
    .clk_2_N_in(clk_2_wires[75]),
    .prog_clk_2_S_out(prog_clk_2_wires[76]),
    .prog_clk_2_N_in(prog_clk_2_wires[75]),
    .prog_clk_0_S_out(prog_clk_0_wires[334]),
    .prog_clk_0_W_in(prog_clk_0_wires[333]),
    .config_enable_S_in(config_enableWires[97]),
    .reset_E_out(resetWires[63]),
    .reset_W_in(resetWires[62]),
    .Test_en_E_out(Test_enWires[63]),
    .Test_en_W_in(Test_enWires[62]),
    .pReset_S_in(pResetWires[97]),
    .chany_bottom_in(sb_1__1__56_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_91_ccff_tail),
    .chany_bottom_out(cby_1__1__81_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__81_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__81_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__81_ccff_tail)
  );


  cby_1__1_
  cby_9__4_
  (
    .clk_2_S_out(clk_2_wires[89]),
    .clk_2_N_in(clk_2_wires[88]),
    .prog_clk_2_S_out(prog_clk_2_wires[89]),
    .prog_clk_2_N_in(prog_clk_2_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[340]),
    .prog_clk_0_W_in(prog_clk_0_wires[339]),
    .config_enable_S_in(config_enableWires[195]),
    .reset_E_out(resetWires[107]),
    .reset_W_in(resetWires[106]),
    .Test_en_E_out(Test_enWires[107]),
    .Test_en_W_in(Test_enWires[106]),
    .pReset_S_in(pResetWires[195]),
    .chany_bottom_in(sb_1__3__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__57_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_92_ccff_tail),
    .chany_bottom_out(cby_1__1__82_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__82_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__82_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__82_ccff_tail)
  );


  cby_1__1_
  cby_9__5_
  (
    .clk_2_N_out(clk_2_wires[87]),
    .clk_2_S_in(clk_2_wires[86]),
    .prog_clk_2_N_out(prog_clk_2_wires[87]),
    .prog_clk_2_S_in(prog_clk_2_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[343]),
    .prog_clk_0_W_in(prog_clk_0_wires[342]),
    .config_enable_S_in(config_enableWires[244]),
    .reset_E_out(resetWires[129]),
    .reset_W_in(resetWires[128]),
    .Test_en_E_out(Test_enWires[129]),
    .Test_en_W_in(Test_enWires[128]),
    .pReset_S_in(pResetWires[244]),
    .chany_bottom_in(sb_1__1__57_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__58_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_93_ccff_tail),
    .chany_bottom_out(cby_1__1__83_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__83_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__83_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__83_ccff_tail)
  );


  cby_1__1_
  cby_9__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[346]),
    .prog_clk_0_W_in(prog_clk_0_wires[345]),
    .config_enable_S_in(config_enableWires[293]),
    .reset_E_out(resetWires[151]),
    .reset_W_in(resetWires[150]),
    .Test_en_E_out(Test_enWires[151]),
    .Test_en_W_in(Test_enWires[150]),
    .pReset_S_in(pResetWires[293]),
    .chany_bottom_in(sb_1__1__58_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__59_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_94_ccff_tail),
    .chany_bottom_out(cby_1__1__84_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__84_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__84_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__84_ccff_tail)
  );


  cby_1__1_
  cby_9__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[349]),
    .prog_clk_0_W_in(prog_clk_0_wires[348]),
    .config_enable_S_in(config_enableWires[342]),
    .reset_E_out(resetWires[173]),
    .reset_W_in(resetWires[172]),
    .Test_en_E_out(Test_enWires[173]),
    .Test_en_W_in(Test_enWires[172]),
    .pReset_S_in(pResetWires[342]),
    .chany_bottom_in(sb_1__1__59_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__60_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_95_ccff_tail),
    .chany_bottom_out(cby_1__1__85_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__85_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__85_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__85_ccff_tail)
  );


  cby_1__1_
  cby_9__8_
  (
    .clk_2_S_out(clk_2_wires[102]),
    .clk_2_N_in(clk_2_wires[101]),
    .prog_clk_2_S_out(prog_clk_2_wires[102]),
    .prog_clk_2_N_in(prog_clk_2_wires[101]),
    .prog_clk_0_S_out(prog_clk_0_wires[352]),
    .prog_clk_0_W_in(prog_clk_0_wires[351]),
    .config_enable_S_in(config_enableWires[391]),
    .reset_E_out(resetWires[195]),
    .reset_W_in(resetWires[194]),
    .Test_en_E_out(Test_enWires[195]),
    .Test_en_W_in(Test_enWires[194]),
    .pReset_S_in(pResetWires[391]),
    .chany_bottom_in(sb_1__1__60_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__61_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_96_ccff_tail),
    .chany_bottom_out(cby_1__1__86_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__86_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__86_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__86_ccff_tail)
  );


  cby_1__1_
  cby_9__9_
  (
    .clk_2_N_out(clk_2_wires[100]),
    .clk_2_S_in(clk_2_wires[99]),
    .prog_clk_2_N_out(prog_clk_2_wires[100]),
    .prog_clk_2_S_in(prog_clk_2_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[355]),
    .prog_clk_0_W_in(prog_clk_0_wires[354]),
    .config_enable_S_in(config_enableWires[440]),
    .reset_E_out(resetWires[217]),
    .reset_W_in(resetWires[216]),
    .Test_en_E_out(Test_enWires[217]),
    .Test_en_W_in(Test_enWires[216]),
    .pReset_S_in(pResetWires[440]),
    .chany_bottom_in(sb_1__1__61_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_97_ccff_tail),
    .chany_bottom_out(cby_1__1__87_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__87_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__87_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__87_ccff_tail)
  );


  cby_1__1_
  cby_9__11_
  (
    .clk_2_N_out(clk_2_wires[111]),
    .clk_2_S_in(clk_2_wires[110]),
    .prog_clk_2_N_out(prog_clk_2_wires[111]),
    .prog_clk_2_S_in(prog_clk_2_wires[110]),
    .prog_clk_0_S_out(prog_clk_0_wires[361]),
    .prog_clk_0_W_in(prog_clk_0_wires[360]),
    .config_enable_S_in(config_enableWires[538]),
    .reset_E_out(resetWires[261]),
    .reset_W_in(resetWires[260]),
    .Test_en_E_out(Test_enWires[261]),
    .Test_en_W_in(Test_enWires[260]),
    .pReset_S_in(pResetWires[538]),
    .chany_bottom_in(sb_1__3__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__62_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_98_ccff_tail),
    .chany_bottom_out(cby_1__1__88_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__88_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__88_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__88_ccff_tail)
  );


  cby_1__1_
  cby_9__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[366]),
    .prog_clk_0_S_out(prog_clk_0_wires[364]),
    .prog_clk_0_W_in(prog_clk_0_wires[363]),
    .config_enable_S_in(config_enableWires[587]),
    .reset_E_out(resetWires[283]),
    .reset_W_in(resetWires[282]),
    .Test_en_E_out(Test_enWires[283]),
    .Test_en_W_in(Test_enWires[282]),
    .pReset_S_in(pResetWires[587]),
    .chany_bottom_in(sb_1__1__62_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__8_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__8_ccff_tail),
    .chany_bottom_out(cby_1__1__89_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__89_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__89_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__89_ccff_tail)
  );


  cby_1__1_
  cby_10__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[369]),
    .prog_clk_0_W_in(prog_clk_0_wires[368]),
    .config_enable_S_in(config_enableWires[54]),
    .reset_E_out(resetWires[43]),
    .reset_W_in(resetWires[42]),
    .Test_en_E_out(Test_enWires[43]),
    .Test_en_W_in(Test_enWires[42]),
    .pReset_S_in(pResetWires[54]),
    .chany_bottom_in(sb_1__0__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__63_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_100_ccff_tail),
    .chany_bottom_out(cby_1__1__90_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__90_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__90_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__90_ccff_tail)
  );


  cby_1__1_
  cby_10__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[372]),
    .prog_clk_0_W_in(prog_clk_0_wires[371]),
    .config_enable_S_in(config_enableWires[101]),
    .reset_E_out(resetWires[65]),
    .reset_W_in(resetWires[64]),
    .Test_en_E_out(Test_enWires[65]),
    .Test_en_W_in(Test_enWires[64]),
    .pReset_S_in(pResetWires[101]),
    .chany_bottom_in(sb_1__1__63_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_101_ccff_tail),
    .chany_bottom_out(cby_1__1__91_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__91_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__91_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__91_ccff_tail)
  );


  cby_1__1_
  cby_10__4_
  (
    .clk_3_S_out(clk_3_wires[83]),
    .clk_3_N_in(clk_3_wires[82]),
    .prog_clk_3_S_out(prog_clk_3_wires[83]),
    .prog_clk_3_N_in(prog_clk_3_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[378]),
    .prog_clk_0_W_in(prog_clk_0_wires[377]),
    .config_enable_S_in(config_enableWires[199]),
    .reset_E_out(resetWires[109]),
    .reset_W_in(resetWires[108]),
    .Test_en_E_out(Test_enWires[109]),
    .Test_en_W_in(Test_enWires[108]),
    .pReset_S_in(pResetWires[199]),
    .chany_bottom_in(sb_2__3__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__64_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_102_ccff_tail),
    .chany_bottom_out(cby_1__1__92_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__92_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__92_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__92_ccff_tail)
  );


  cby_1__1_
  cby_10__5_
  (
    .clk_3_S_out(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[76]),
    .prog_clk_3_S_out(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[381]),
    .prog_clk_0_W_in(prog_clk_0_wires[380]),
    .config_enable_S_in(config_enableWires[248]),
    .reset_E_out(resetWires[131]),
    .reset_W_in(resetWires[130]),
    .Test_en_E_out(Test_enWires[131]),
    .Test_en_W_in(Test_enWires[130]),
    .pReset_S_in(pResetWires[248]),
    .chany_bottom_in(sb_1__1__64_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__65_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_103_ccff_tail),
    .chany_bottom_out(cby_1__1__93_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__93_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__93_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__93_ccff_tail)
  );


  cby_1__1_
  cby_10__6_
  (
    .clk_3_S_out(clk_3_wires[73]),
    .clk_3_N_in(clk_3_wires[72]),
    .prog_clk_3_S_out(prog_clk_3_wires[73]),
    .prog_clk_3_N_in(prog_clk_3_wires[72]),
    .prog_clk_0_S_out(prog_clk_0_wires[384]),
    .prog_clk_0_W_in(prog_clk_0_wires[383]),
    .config_enable_S_in(config_enableWires[297]),
    .reset_E_out(resetWires[153]),
    .reset_W_in(resetWires[152]),
    .Test_en_E_out(Test_enWires[153]),
    .Test_en_W_in(Test_enWires[152]),
    .pReset_S_in(pResetWires[297]),
    .chany_bottom_in(sb_1__1__65_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__66_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_104_ccff_tail),
    .chany_bottom_out(cby_1__1__94_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__94_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__94_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__94_ccff_tail)
  );


  cby_1__1_
  cby_10__7_
  (
    .clk_3_N_out(clk_3_wires[71]),
    .clk_3_S_in(clk_3_wires[70]),
    .prog_clk_3_N_out(prog_clk_3_wires[71]),
    .prog_clk_3_S_in(prog_clk_3_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[387]),
    .prog_clk_0_W_in(prog_clk_0_wires[386]),
    .config_enable_S_in(config_enableWires[346]),
    .reset_E_out(resetWires[175]),
    .reset_W_in(resetWires[174]),
    .Test_en_E_out(Test_enWires[175]),
    .Test_en_W_in(Test_enWires[174]),
    .pReset_S_in(pResetWires[346]),
    .chany_bottom_in(sb_1__1__66_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__67_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_105_ccff_tail),
    .chany_bottom_out(cby_1__1__95_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__95_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__95_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__95_ccff_tail)
  );


  cby_1__1_
  cby_10__8_
  (
    .clk_3_N_out(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[74]),
    .prog_clk_3_N_out(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[74]),
    .prog_clk_0_S_out(prog_clk_0_wires[390]),
    .prog_clk_0_W_in(prog_clk_0_wires[389]),
    .config_enable_S_in(config_enableWires[395]),
    .reset_E_out(resetWires[197]),
    .reset_W_in(resetWires[196]),
    .Test_en_E_out(Test_enWires[197]),
    .Test_en_W_in(Test_enWires[196]),
    .pReset_S_in(pResetWires[395]),
    .chany_bottom_in(sb_1__1__67_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__68_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_106_ccff_tail),
    .chany_bottom_out(cby_1__1__96_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__96_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__96_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__96_ccff_tail)
  );


  cby_1__1_
  cby_10__9_
  (
    .clk_3_N_out(clk_3_wires[81]),
    .clk_3_S_in(clk_3_wires[80]),
    .prog_clk_3_N_out(prog_clk_3_wires[81]),
    .prog_clk_3_S_in(prog_clk_3_wires[80]),
    .prog_clk_0_S_out(prog_clk_0_wires[393]),
    .prog_clk_0_W_in(prog_clk_0_wires[392]),
    .config_enable_S_in(config_enableWires[444]),
    .reset_E_out(resetWires[219]),
    .reset_W_in(resetWires[218]),
    .Test_en_E_out(Test_enWires[219]),
    .Test_en_W_in(Test_enWires[218]),
    .pReset_S_in(pResetWires[444]),
    .chany_bottom_in(sb_1__1__68_chany_top_out[0:19]),
    .chany_top_in(sb_2__2__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_107_ccff_tail),
    .chany_bottom_out(cby_1__1__97_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__97_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__97_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__97_ccff_tail)
  );


  cby_1__1_
  cby_10__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[399]),
    .prog_clk_0_W_in(prog_clk_0_wires[398]),
    .config_enable_S_in(config_enableWires[542]),
    .reset_E_out(resetWires[263]),
    .reset_W_in(resetWires[262]),
    .Test_en_E_out(Test_enWires[263]),
    .Test_en_W_in(Test_enWires[262]),
    .pReset_S_in(pResetWires[542]),
    .chany_bottom_in(sb_2__3__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__69_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_108_ccff_tail),
    .chany_bottom_out(cby_1__1__98_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__98_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__98_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__98_ccff_tail)
  );


  cby_1__1_
  cby_10__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[404]),
    .prog_clk_0_S_out(prog_clk_0_wires[402]),
    .prog_clk_0_W_in(prog_clk_0_wires[401]),
    .config_enable_S_in(config_enableWires[591]),
    .reset_E_out(resetWires[285]),
    .reset_W_in(resetWires[284]),
    .Test_en_E_out(Test_enWires[285]),
    .Test_en_W_in(Test_enWires[284]),
    .pReset_S_in(pResetWires[591]),
    .chany_bottom_in(sb_1__1__69_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__9_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__9_ccff_tail),
    .chany_bottom_out(cby_1__1__99_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__99_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__99_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__99_ccff_tail)
  );


  cby_1__1_
  cby_11__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[407]),
    .prog_clk_0_W_in(prog_clk_0_wires[406]),
    .config_enable_S_in(config_enableWires[57]),
    .reset_E_out(resetWires[45]),
    .reset_W_in(resetWires[44]),
    .Test_en_E_out(Test_enWires[45]),
    .Test_en_W_in(Test_enWires[44]),
    .pReset_S_in(pResetWires[57]),
    .chany_bottom_in(sb_1__0__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__70_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_110_ccff_tail),
    .chany_bottom_out(cby_1__1__100_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__100_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__100_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__100_ccff_tail)
  );


  cby_1__1_
  cby_11__2_
  (
    .clk_2_S_out(clk_2_wires[116]),
    .clk_2_N_in(clk_2_wires[115]),
    .prog_clk_2_S_out(prog_clk_2_wires[116]),
    .prog_clk_2_N_in(prog_clk_2_wires[115]),
    .prog_clk_0_S_out(prog_clk_0_wires[410]),
    .prog_clk_0_W_in(prog_clk_0_wires[409]),
    .config_enable_S_in(config_enableWires[105]),
    .reset_E_out(resetWires[67]),
    .reset_W_in(resetWires[66]),
    .Test_en_E_out(Test_enWires[67]),
    .Test_en_W_in(Test_enWires[66]),
    .pReset_S_in(pResetWires[105]),
    .chany_bottom_in(sb_1__1__70_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_111_ccff_tail),
    .chany_bottom_out(cby_1__1__101_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__101_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__101_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__101_ccff_tail)
  );


  cby_1__1_
  cby_11__4_
  (
    .clk_2_S_out(clk_2_wires[123]),
    .clk_2_N_in(clk_2_wires[122]),
    .prog_clk_2_S_out(prog_clk_2_wires[123]),
    .prog_clk_2_N_in(prog_clk_2_wires[122]),
    .prog_clk_0_S_out(prog_clk_0_wires[416]),
    .prog_clk_0_W_in(prog_clk_0_wires[415]),
    .config_enable_S_in(config_enableWires[203]),
    .reset_E_out(resetWires[111]),
    .reset_W_in(resetWires[110]),
    .Test_en_E_out(Test_enWires[111]),
    .Test_en_W_in(Test_enWires[110]),
    .pReset_S_in(pResetWires[203]),
    .chany_bottom_in(sb_1__3__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__71_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_112_ccff_tail),
    .chany_bottom_out(cby_1__1__102_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__102_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__102_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__102_ccff_tail)
  );


  cby_1__1_
  cby_11__5_
  (
    .clk_2_N_out(clk_2_wires[121]),
    .clk_2_S_in(clk_2_wires[120]),
    .prog_clk_2_N_out(prog_clk_2_wires[121]),
    .prog_clk_2_S_in(prog_clk_2_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[419]),
    .prog_clk_0_W_in(prog_clk_0_wires[418]),
    .config_enable_S_in(config_enableWires[252]),
    .reset_E_out(resetWires[133]),
    .reset_W_in(resetWires[132]),
    .Test_en_E_out(Test_enWires[133]),
    .Test_en_W_in(Test_enWires[132]),
    .pReset_S_in(pResetWires[252]),
    .chany_bottom_in(sb_1__1__71_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__72_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_113_ccff_tail),
    .chany_bottom_out(cby_1__1__103_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__103_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__103_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__103_ccff_tail)
  );


  cby_1__1_
  cby_11__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[422]),
    .prog_clk_0_W_in(prog_clk_0_wires[421]),
    .config_enable_S_in(config_enableWires[301]),
    .reset_E_out(resetWires[155]),
    .reset_W_in(resetWires[154]),
    .Test_en_E_out(Test_enWires[155]),
    .Test_en_W_in(Test_enWires[154]),
    .pReset_S_in(pResetWires[301]),
    .chany_bottom_in(sb_1__1__72_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__73_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_114_ccff_tail),
    .chany_bottom_out(cby_1__1__104_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__104_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__104_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__104_ccff_tail)
  );


  cby_1__1_
  cby_11__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[425]),
    .prog_clk_0_W_in(prog_clk_0_wires[424]),
    .config_enable_S_in(config_enableWires[350]),
    .reset_E_out(resetWires[177]),
    .reset_W_in(resetWires[176]),
    .Test_en_E_out(Test_enWires[177]),
    .Test_en_W_in(Test_enWires[176]),
    .pReset_S_in(pResetWires[350]),
    .chany_bottom_in(sb_1__1__73_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__74_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_115_ccff_tail),
    .chany_bottom_out(cby_1__1__105_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__105_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__105_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__105_ccff_tail)
  );


  cby_1__1_
  cby_11__8_
  (
    .clk_2_S_out(clk_2_wires[130]),
    .clk_2_N_in(clk_2_wires[129]),
    .prog_clk_2_S_out(prog_clk_2_wires[130]),
    .prog_clk_2_N_in(prog_clk_2_wires[129]),
    .prog_clk_0_S_out(prog_clk_0_wires[428]),
    .prog_clk_0_W_in(prog_clk_0_wires[427]),
    .config_enable_S_in(config_enableWires[399]),
    .reset_E_out(resetWires[199]),
    .reset_W_in(resetWires[198]),
    .Test_en_E_out(Test_enWires[199]),
    .Test_en_W_in(Test_enWires[198]),
    .pReset_S_in(pResetWires[399]),
    .chany_bottom_in(sb_1__1__74_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__75_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_116_ccff_tail),
    .chany_bottom_out(cby_1__1__106_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__106_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__106_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__106_ccff_tail)
  );


  cby_1__1_
  cby_11__9_
  (
    .clk_2_N_out(clk_2_wires[128]),
    .clk_2_S_in(clk_2_wires[127]),
    .prog_clk_2_N_out(prog_clk_2_wires[128]),
    .prog_clk_2_S_in(prog_clk_2_wires[127]),
    .prog_clk_0_S_out(prog_clk_0_wires[431]),
    .prog_clk_0_W_in(prog_clk_0_wires[430]),
    .config_enable_S_in(config_enableWires[448]),
    .reset_E_out(resetWires[221]),
    .reset_W_in(resetWires[220]),
    .Test_en_E_out(Test_enWires[221]),
    .Test_en_W_in(Test_enWires[220]),
    .pReset_S_in(pResetWires[448]),
    .chany_bottom_in(sb_1__1__75_chany_top_out[0:19]),
    .chany_top_in(sb_1__2__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_117_ccff_tail),
    .chany_bottom_out(cby_1__1__107_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__107_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__107_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__107_ccff_tail)
  );


  cby_1__1_
  cby_11__11_
  (
    .clk_2_N_out(clk_2_wires[135]),
    .clk_2_S_in(clk_2_wires[134]),
    .prog_clk_2_N_out(prog_clk_2_wires[135]),
    .prog_clk_2_S_in(prog_clk_2_wires[134]),
    .prog_clk_0_S_out(prog_clk_0_wires[437]),
    .prog_clk_0_W_in(prog_clk_0_wires[436]),
    .config_enable_S_in(config_enableWires[546]),
    .reset_E_out(resetWires[265]),
    .reset_W_in(resetWires[264]),
    .Test_en_E_out(Test_enWires[265]),
    .Test_en_W_in(Test_enWires[264]),
    .pReset_S_in(pResetWires[546]),
    .chany_bottom_in(sb_1__3__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__76_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_118_ccff_tail),
    .chany_bottom_out(cby_1__1__108_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__108_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__108_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__108_ccff_tail)
  );


  cby_1__1_
  cby_11__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[442]),
    .prog_clk_0_S_out(prog_clk_0_wires[440]),
    .prog_clk_0_W_in(prog_clk_0_wires[439]),
    .config_enable_S_in(config_enableWires[595]),
    .reset_E_out(resetWires[287]),
    .reset_W_in(resetWires[286]),
    .Test_en_E_out(Test_enWires[287]),
    .Test_en_W_in(Test_enWires[286]),
    .pReset_S_in(pResetWires[595]),
    .chany_bottom_in(sb_1__1__76_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__10_chany_bottom_out[0:19]),
    .ccff_head(sb_1__12__10_ccff_tail),
    .chany_bottom_out(cby_1__1__109_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__109_chany_top_out[0:19]),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
    .left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__109_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
    .ccff_tail(cby_1__1__109_ccff_tail)
  );


  cby_2__3_
  cby_2__3_
  (
    .clk_3_S_out(clk_3_wires[69]),
    .clk_3_N_in(clk_3_wires[68]),
    .prog_clk_3_S_out(prog_clk_3_wires[69]),
    .prog_clk_3_N_in(prog_clk_3_wires[68]),
    .prog_clk_0_S_out(prog_clk_0_wires[71]),
    .prog_clk_0_W_in(prog_clk_0_wires[70]),
    .config_enable_S_in(config_enableWires[118]),
    .reset_E_in(resetWires[72]),
    .reset_W_out(resetWires[69]),
    .Test_en_E_in(Test_enWires[72]),
    .Test_en_W_out(Test_enWires[69]),
    .pReset_S_in(pResetWires[118]),
    .chany_bottom_in(sb_2__2__0_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__0_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_2_ccff_tail),
    .chany_bottom_out(cby_2__3__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__0_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__0_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__0_ccff_tail)
  );


  cby_2__3_
  cby_2__10_
  (
    .clk_3_N_out(clk_3_wires[67]),
    .clk_3_S_in(clk_3_wires[66]),
    .prog_clk_3_N_out(prog_clk_3_wires[67]),
    .prog_clk_3_S_in(prog_clk_3_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[92]),
    .prog_clk_0_W_in(prog_clk_0_wires[91]),
    .config_enable_S_in(config_enableWires[461]),
    .reset_E_in(resetWires[226]),
    .reset_W_out(resetWires[223]),
    .Test_en_E_in(Test_enWires[226]),
    .Test_en_W_out(Test_enWires[223]),
    .pReset_S_in(pResetWires[461]),
    .chany_bottom_in(sb_2__2__1_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__1_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_3_ccff_tail),
    .chany_bottom_out(cby_2__3__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__1_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__1_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__1_ccff_tail)
  );


  cby_2__3_
  cby_4__3_
  (
    .clk_3_S_out(clk_3_wires[25]),
    .clk_3_N_in(clk_3_wires[24]),
    .prog_clk_3_S_out(prog_clk_3_wires[25]),
    .prog_clk_3_N_in(prog_clk_3_wires[24]),
    .prog_clk_0_S_out(prog_clk_0_wires[147]),
    .prog_clk_0_W_in(prog_clk_0_wires[146]),
    .config_enable_S_in(config_enableWires[126]),
    .reset_E_in(resetWires[76]),
    .reset_W_out(resetWires[73]),
    .Test_en_E_in(Test_enWires[76]),
    .Test_en_W_out(Test_enWires[73]),
    .pReset_S_in(pResetWires[126]),
    .chany_bottom_in(sb_2__2__2_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__2_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_4_ccff_tail),
    .chany_bottom_out(cby_2__3__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__2_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__2_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__2_ccff_tail)
  );


  cby_2__3_
  cby_4__10_
  (
    .clk_3_N_out(clk_3_wires[23]),
    .clk_3_S_in(clk_3_wires[22]),
    .prog_clk_3_N_out(prog_clk_3_wires[23]),
    .prog_clk_3_S_in(prog_clk_3_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[168]),
    .prog_clk_0_W_in(prog_clk_0_wires[167]),
    .config_enable_S_in(config_enableWires[469]),
    .reset_E_in(resetWires[230]),
    .reset_W_out(resetWires[227]),
    .Test_en_E_in(Test_enWires[230]),
    .Test_en_W_out(Test_enWires[227]),
    .pReset_S_in(pResetWires[469]),
    .chany_bottom_in(sb_2__2__3_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__3_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_5_ccff_tail),
    .chany_bottom_out(cby_2__3__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__3_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__3_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__3_ccff_tail)
  );


  cby_2__3_
  cby_6__3_
  (
    .clk_3_S_in(clk_3_wires[94]),
    .clk_3_N_out(clk_3_wires[93]),
    .prog_clk_3_S_in(prog_clk_3_wires[94]),
    .prog_clk_3_N_out(prog_clk_3_wires[93]),
    .prog_clk_0_S_out(prog_clk_0_wires[223]),
    .prog_clk_0_W_in(prog_clk_0_wires[222]),
    .config_enable_N_out(config_enableWires[6]),
    .config_enable_S_in(config_enableWires[134]),
    .reset_E_out(resetWires[79]),
    .reset_W_out(resetWires[77]),
    .reset_N_out(resetWires[6]),
    .reset_S_in(resetWires[5]),
    .Test_en_E_out(Test_enWires[79]),
    .Test_en_W_out(Test_enWires[77]),
    .Test_en_N_out(Test_enWires[6]),
    .Test_en_S_in(Test_enWires[5]),
    .pReset_N_out(pResetWires[6]),
    .pReset_S_in(pResetWires[134]),
    .chany_bottom_in(sb_2__2__4_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__4_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_6_ccff_tail),
    .chany_bottom_out(cby_2__3__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__4_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__4_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__4_ccff_tail)
  );


  cby_2__3_
  cby_6__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[244]),
    .prog_clk_0_W_in(prog_clk_0_wires[243]),
    .config_enable_N_out(config_enableWires[20]),
    .config_enable_S_in(config_enableWires[477]),
    .reset_E_out(resetWires[233]),
    .reset_W_out(resetWires[231]),
    .reset_N_out(resetWires[20]),
    .reset_S_in(resetWires[19]),
    .Test_en_E_out(Test_enWires[233]),
    .Test_en_W_out(Test_enWires[231]),
    .Test_en_N_out(Test_enWires[20]),
    .Test_en_S_in(Test_enWires[19]),
    .pReset_N_out(pResetWires[20]),
    .pReset_S_in(pResetWires[477]),
    .chany_bottom_in(sb_2__2__5_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__5_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_7_ccff_tail),
    .chany_bottom_out(cby_2__3__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__5_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__5_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__5_ccff_tail)
  );


  cby_2__3_
  cby_8__3_
  (
    .clk_3_S_out(clk_3_wires[43]),
    .clk_3_N_in(clk_3_wires[42]),
    .prog_clk_3_S_out(prog_clk_3_wires[43]),
    .prog_clk_3_N_in(prog_clk_3_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[299]),
    .prog_clk_0_W_in(prog_clk_0_wires[298]),
    .config_enable_S_in(config_enableWires[142]),
    .reset_E_out(resetWires[83]),
    .reset_W_in(resetWires[82]),
    .Test_en_E_out(Test_enWires[83]),
    .Test_en_W_in(Test_enWires[82]),
    .pReset_S_in(pResetWires[142]),
    .chany_bottom_in(sb_2__2__6_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__6_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_8_ccff_tail),
    .chany_bottom_out(cby_2__3__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__6_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__6_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__6_ccff_tail)
  );


  cby_2__3_
  cby_8__10_
  (
    .clk_3_N_out(clk_3_wires[41]),
    .clk_3_S_in(clk_3_wires[40]),
    .prog_clk_3_N_out(prog_clk_3_wires[41]),
    .prog_clk_3_S_in(prog_clk_3_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[320]),
    .prog_clk_0_W_in(prog_clk_0_wires[319]),
    .config_enable_S_in(config_enableWires[485]),
    .reset_E_out(resetWires[237]),
    .reset_W_in(resetWires[236]),
    .Test_en_E_out(Test_enWires[237]),
    .Test_en_W_in(Test_enWires[236]),
    .pReset_S_in(pResetWires[485]),
    .chany_bottom_in(sb_2__2__7_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__7_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_9_ccff_tail),
    .chany_bottom_out(cby_2__3__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__7_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__7_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__7_ccff_tail)
  );


  cby_2__3_
  cby_10__3_
  (
    .clk_3_S_out(clk_3_wires[87]),
    .clk_3_N_in(clk_3_wires[86]),
    .prog_clk_3_S_out(prog_clk_3_wires[87]),
    .prog_clk_3_N_in(prog_clk_3_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[375]),
    .prog_clk_0_W_in(prog_clk_0_wires[374]),
    .config_enable_S_in(config_enableWires[150]),
    .reset_E_out(resetWires[87]),
    .reset_W_in(resetWires[86]),
    .Test_en_E_out(Test_enWires[87]),
    .Test_en_W_in(Test_enWires[86]),
    .pReset_S_in(pResetWires[150]),
    .chany_bottom_in(sb_2__2__8_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__8_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_10_ccff_tail),
    .chany_bottom_out(cby_2__3__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__8_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__8_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__8_ccff_tail)
  );


  cby_2__3_
  cby_10__10_
  (
    .clk_3_N_out(clk_3_wires[85]),
    .clk_3_S_in(clk_3_wires[84]),
    .prog_clk_3_N_out(prog_clk_3_wires[85]),
    .prog_clk_3_S_in(prog_clk_3_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[396]),
    .prog_clk_0_W_in(prog_clk_0_wires[395]),
    .config_enable_S_in(config_enableWires[493]),
    .reset_E_out(resetWires[241]),
    .reset_W_in(resetWires[240]),
    .Test_en_E_out(Test_enWires[241]),
    .Test_en_W_in(Test_enWires[240]),
    .pReset_S_in(pResetWires[493]),
    .chany_bottom_in(sb_2__2__9_chany_top_out[0:19]),
    .chany_top_in(sb_2__3__9_chany_bottom_out[0:19]),
    .ccff_head(grid_mult_18_11_ccff_tail),
    .chany_bottom_out(cby_2__3__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_2__3__9_chany_top_out[0:19]),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_a_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_a_17_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_12_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_12_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_13_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_13_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_14_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_14_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_15_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_15_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_16_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_16_),
    .left_grid_right_width_1_height_0_subtile_0__pin_b_17_(cby_2__3__9_left_grid_right_width_1_height_0_subtile_0__pin_b_17_),
    .ccff_tail(cby_2__3__9_ccff_tail)
  );


  cby_4__1_
  cby_12__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[445]),
    .prog_clk_0_W_in(prog_clk_0_wires[444]),
    .config_enable_S_in(config_enableWires[60]),
    .pReset_S_in(pResetWires[60]),
    .chany_bottom_in(sb_12__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[11]),
    .chany_bottom_out(cby_12__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__0_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[23]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[23]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[23]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_11_ccff_tail)
  );


  cby_4__1_
  cby_12__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[448]),
    .prog_clk_0_W_in(prog_clk_0_wires[447]),
    .config_enable_S_in(config_enableWires[109]),
    .pReset_S_in(pResetWires[109]),
    .chany_bottom_in(sb_12__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__2__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[10]),
    .chany_bottom_out(cby_12__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__1_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[22]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[22]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[22]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_10_ccff_tail)
  );


  cby_4__1_
  cby_12__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[454]),
    .prog_clk_0_W_in(prog_clk_0_wires[453]),
    .config_enable_S_in(config_enableWires[207]),
    .pReset_S_in(pResetWires[207]),
    .chany_bottom_in(sb_12__3__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[8]),
    .chany_bottom_out(cby_12__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__2_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[20]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[20]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[20]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_8_ccff_tail)
  );


  cby_4__1_
  cby_12__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[457]),
    .prog_clk_0_W_in(prog_clk_0_wires[456]),
    .config_enable_S_in(config_enableWires[256]),
    .pReset_S_in(pResetWires[256]),
    .chany_bottom_in(sb_12__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__2_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[7]),
    .chany_bottom_out(cby_12__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__3_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[19]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[19]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[19]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_7_ccff_tail)
  );


  cby_4__1_
  cby_12__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[460]),
    .prog_clk_0_W_in(prog_clk_0_wires[459]),
    .config_enable_S_in(config_enableWires[305]),
    .pReset_S_in(pResetWires[305]),
    .chany_bottom_in(sb_12__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__3_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[6]),
    .chany_bottom_out(cby_12__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__4_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[18]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[18]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[18]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_6_ccff_tail)
  );


  cby_4__1_
  cby_12__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[463]),
    .prog_clk_0_W_in(prog_clk_0_wires[462]),
    .config_enable_S_in(config_enableWires[354]),
    .pReset_S_in(pResetWires[354]),
    .chany_bottom_in(sb_12__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__4_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[5]),
    .chany_bottom_out(cby_12__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__5_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[17]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[17]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[17]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_5_ccff_tail)
  );


  cby_4__1_
  cby_12__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[466]),
    .prog_clk_0_W_in(prog_clk_0_wires[465]),
    .config_enable_S_in(config_enableWires[403]),
    .pReset_S_in(pResetWires[403]),
    .chany_bottom_in(sb_12__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__5_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[4]),
    .chany_bottom_out(cby_12__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__6_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[16]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[16]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[16]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_4_ccff_tail)
  );


  cby_4__1_
  cby_12__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[469]),
    .prog_clk_0_W_in(prog_clk_0_wires[468]),
    .config_enable_S_in(config_enableWires[452]),
    .pReset_S_in(pResetWires[452]),
    .chany_bottom_in(sb_12__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_12__2__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[3]),
    .chany_bottom_out(cby_12__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__7_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[15]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[15]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[15]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_3_ccff_tail)
  );


  cby_4__1_
  cby_12__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[475]),
    .prog_clk_0_W_in(prog_clk_0_wires[474]),
    .config_enable_S_in(config_enableWires[550]),
    .pReset_S_in(pResetWires[550]),
    .chany_bottom_in(sb_12__3__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__6_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[1]),
    .chany_bottom_out(cby_12__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__8_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[13]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[13]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[13]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_1_ccff_tail)
  );


  cby_4__1_
  cby_12__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[480]),
    .prog_clk_0_S_out(prog_clk_0_wires[478]),
    .prog_clk_0_W_in(prog_clk_0_wires[477]),
    .config_enable_S_in(config_enableWires[599]),
    .pReset_S_in(pResetWires[599]),
    .chany_bottom_in(sb_12__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_12__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_12__12__0_ccff_tail),
    .chany_bottom_out(cby_12__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__9_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[12]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[12]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[12]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_0_ccff_tail)
  );


  cby_4__3_
  cby_12__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[451]),
    .prog_clk_0_W_in(prog_clk_0_wires[450]),
    .config_enable_S_in(config_enableWires[158]),
    .pReset_S_in(pResetWires[158]),
    .chany_bottom_in(sb_12__2__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__3__0_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[9]),
    .chany_bottom_out(cby_12__3__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__3__0_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[21]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[21]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[21]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_9_ccff_tail)
  );


  cby_4__3_
  cby_12__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[472]),
    .prog_clk_0_W_in(prog_clk_0_wires[471]),
    .config_enable_S_in(config_enableWires[501]),
    .pReset_S_in(pResetWires[501]),
    .chany_bottom_in(sb_12__2__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__3__1_chany_bottom_out[0:19]),
    .ccff_head(ccff_head[2]),
    .chany_bottom_out(cby_12__3__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__3__1_chany_top_out[0:19]),
    .IO_ISOL_N(IO_ISOL_N),
    .gfpga_pad_sofa_plus_io_SOC_IN(gfpga_pad_sofa_plus_io_SOC_IN[14]),
    .gfpga_pad_sofa_plus_io_SOC_OUT(gfpga_pad_sofa_plus_io_SOC_OUT[14]),
    .gfpga_pad_sofa_plus_io_SOC_DIR(gfpga_pad_sofa_plus_io_SOC_DIR[14]),
    .left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
    .left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
    .ccff_tail(grid_io_right_right_2_ccff_tail)
  );


  direct_interc
  direct_interc_0_
  (
    .in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_0_out)
  );


  direct_interc
  direct_interc_1_
  (
    .in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_1_out)
  );


  direct_interc
  direct_interc_2_
  (
    .in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_2_out)
  );


  direct_interc
  direct_interc_3_
  (
    .in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_3_out)
  );


  direct_interc
  direct_interc_4_
  (
    .in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_4_out)
  );


  direct_interc
  direct_interc_5_
  (
    .in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_5_out)
  );


  direct_interc
  direct_interc_6_
  (
    .in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_6_out)
  );


  direct_interc
  direct_interc_7_
  (
    .in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_7_out)
  );


  direct_interc
  direct_interc_8_
  (
    .in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_8_out)
  );


  direct_interc
  direct_interc_9_
  (
    .in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_9_out)
  );


  direct_interc
  direct_interc_10_
  (
    .in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_10_out)
  );


  direct_interc
  direct_interc_11_
  (
    .in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_11_out)
  );


  direct_interc
  direct_interc_12_
  (
    .in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_12_out)
  );


  direct_interc
  direct_interc_13_
  (
    .in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_13_out)
  );


  direct_interc
  direct_interc_14_
  (
    .in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_14_out)
  );


  direct_interc
  direct_interc_15_
  (
    .in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_15_out)
  );


  direct_interc
  direct_interc_16_
  (
    .in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_16_out)
  );


  direct_interc
  direct_interc_17_
  (
    .in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_17_out)
  );


  direct_interc
  direct_interc_18_
  (
    .in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_18_out)
  );


  direct_interc
  direct_interc_19_
  (
    .in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_19_out)
  );


  direct_interc
  direct_interc_20_
  (
    .in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_20_out)
  );


  direct_interc
  direct_interc_21_
  (
    .in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_21_out)
  );


  direct_interc
  direct_interc_22_
  (
    .in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_22_out)
  );


  direct_interc
  direct_interc_23_
  (
    .in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_23_out)
  );


  direct_interc
  direct_interc_24_
  (
    .in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_24_out)
  );


  direct_interc
  direct_interc_25_
  (
    .in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_25_out)
  );


  direct_interc
  direct_interc_26_
  (
    .in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_26_out)
  );


  direct_interc
  direct_interc_27_
  (
    .in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_27_out)
  );


  direct_interc
  direct_interc_28_
  (
    .in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_28_out)
  );


  direct_interc
  direct_interc_29_
  (
    .in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_29_out)
  );


  direct_interc
  direct_interc_30_
  (
    .in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_30_out)
  );


  direct_interc
  direct_interc_31_
  (
    .in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_31_out)
  );


  direct_interc
  direct_interc_32_
  (
    .in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_32_out)
  );


  direct_interc
  direct_interc_33_
  (
    .in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_33_out)
  );


  direct_interc
  direct_interc_34_
  (
    .in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_34_out)
  );


  direct_interc
  direct_interc_35_
  (
    .in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_35_out)
  );


  direct_interc
  direct_interc_36_
  (
    .in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_36_out)
  );


  direct_interc
  direct_interc_37_
  (
    .in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_37_out)
  );


  direct_interc
  direct_interc_38_
  (
    .in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_38_out)
  );


  direct_interc
  direct_interc_39_
  (
    .in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_39_out)
  );


  direct_interc
  direct_interc_40_
  (
    .in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_40_out)
  );


  direct_interc
  direct_interc_41_
  (
    .in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_41_out)
  );


  direct_interc
  direct_interc_42_
  (
    .in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_42_out)
  );


  direct_interc
  direct_interc_43_
  (
    .in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_43_out)
  );


  direct_interc
  direct_interc_44_
  (
    .in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_44_out)
  );


  direct_interc
  direct_interc_45_
  (
    .in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_45_out)
  );


  direct_interc
  direct_interc_46_
  (
    .in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_46_out)
  );


  direct_interc
  direct_interc_47_
  (
    .in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_47_out)
  );


  direct_interc
  direct_interc_48_
  (
    .in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_48_out)
  );


  direct_interc
  direct_interc_49_
  (
    .in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_49_out)
  );


  direct_interc
  direct_interc_50_
  (
    .in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_50_out)
  );


  direct_interc
  direct_interc_51_
  (
    .in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_51_out)
  );


  direct_interc
  direct_interc_52_
  (
    .in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_52_out)
  );


  direct_interc
  direct_interc_53_
  (
    .in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_53_out)
  );


  direct_interc
  direct_interc_54_
  (
    .in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_54_out)
  );


  direct_interc
  direct_interc_55_
  (
    .in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_55_out)
  );


  direct_interc
  direct_interc_56_
  (
    .in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_56_out)
  );


  direct_interc
  direct_interc_57_
  (
    .in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_57_out)
  );


  direct_interc
  direct_interc_58_
  (
    .in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_58_out)
  );


  direct_interc
  direct_interc_59_
  (
    .in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_59_out)
  );


  direct_interc
  direct_interc_60_
  (
    .in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_60_out)
  );


  direct_interc
  direct_interc_61_
  (
    .in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_61_out)
  );


  direct_interc
  direct_interc_62_
  (
    .in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_62_out)
  );


  direct_interc
  direct_interc_63_
  (
    .in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_63_out)
  );


  direct_interc
  direct_interc_64_
  (
    .in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_64_out)
  );


  direct_interc
  direct_interc_65_
  (
    .in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_65_out)
  );


  direct_interc
  direct_interc_66_
  (
    .in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_66_out)
  );


  direct_interc
  direct_interc_67_
  (
    .in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_67_out)
  );


  direct_interc
  direct_interc_68_
  (
    .in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_68_out)
  );


  direct_interc
  direct_interc_69_
  (
    .in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_69_out)
  );


  direct_interc
  direct_interc_70_
  (
    .in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_70_out)
  );


  direct_interc
  direct_interc_71_
  (
    .in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_71_out)
  );


  direct_interc
  direct_interc_72_
  (
    .in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_72_out)
  );


  direct_interc
  direct_interc_73_
  (
    .in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_73_out)
  );


  direct_interc
  direct_interc_74_
  (
    .in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_74_out)
  );


  direct_interc
  direct_interc_75_
  (
    .in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_75_out)
  );


  direct_interc
  direct_interc_76_
  (
    .in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_76_out)
  );


  direct_interc
  direct_interc_77_
  (
    .in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_77_out)
  );


  direct_interc
  direct_interc_78_
  (
    .in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_78_out)
  );


  direct_interc
  direct_interc_79_
  (
    .in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_79_out)
  );


  direct_interc
  direct_interc_80_
  (
    .in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_80_out)
  );


  direct_interc
  direct_interc_81_
  (
    .in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_81_out)
  );


  direct_interc
  direct_interc_82_
  (
    .in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_82_out)
  );


  direct_interc
  direct_interc_83_
  (
    .in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_cout_0_),
    .out(direct_interc_83_out)
  );


  direct_interc
  direct_interc_84_
  (
    .in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_84_out)
  );


  direct_interc
  direct_interc_85_
  (
    .in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_85_out)
  );


  direct_interc
  direct_interc_86_
  (
    .in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_86_out)
  );


  direct_interc
  direct_interc_87_
  (
    .in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_87_out)
  );


  direct_interc
  direct_interc_88_
  (
    .in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_88_out)
  );


  direct_interc
  direct_interc_89_
  (
    .in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_89_out)
  );


  direct_interc
  direct_interc_90_
  (
    .in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_90_out)
  );


  direct_interc
  direct_interc_91_
  (
    .in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_91_out)
  );


  direct_interc
  direct_interc_92_
  (
    .in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_92_out)
  );


  direct_interc
  direct_interc_93_
  (
    .in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_93_out)
  );


  direct_interc
  direct_interc_94_
  (
    .in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_94_out)
  );


  direct_interc
  direct_interc_95_
  (
    .in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_95_out)
  );


  direct_interc
  direct_interc_96_
  (
    .in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_96_out)
  );


  direct_interc
  direct_interc_97_
  (
    .in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_97_out)
  );


  direct_interc
  direct_interc_98_
  (
    .in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_98_out)
  );


  direct_interc
  direct_interc_99_
  (
    .in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_99_out)
  );


  direct_interc
  direct_interc_100_
  (
    .in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_100_out)
  );


  direct_interc
  direct_interc_101_
  (
    .in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_101_out)
  );


  direct_interc
  direct_interc_102_
  (
    .in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_102_out)
  );


  direct_interc
  direct_interc_103_
  (
    .in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_103_out)
  );


  direct_interc
  direct_interc_104_
  (
    .in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_104_out)
  );


  direct_interc
  direct_interc_105_
  (
    .in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_105_out)
  );


  direct_interc
  direct_interc_106_
  (
    .in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_106_out)
  );


  direct_interc
  direct_interc_107_
  (
    .in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_107_out)
  );


  direct_interc
  direct_interc_108_
  (
    .in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_108_out)
  );


  direct_interc
  direct_interc_109_
  (
    .in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_109_out)
  );


  direct_interc
  direct_interc_110_
  (
    .in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_110_out)
  );


  direct_interc
  direct_interc_111_
  (
    .in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_111_out)
  );


  direct_interc
  direct_interc_112_
  (
    .in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_112_out)
  );


  direct_interc
  direct_interc_113_
  (
    .in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_113_out)
  );


  direct_interc
  direct_interc_114_
  (
    .in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_114_out)
  );


  direct_interc
  direct_interc_115_
  (
    .in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_115_out)
  );


  direct_interc
  direct_interc_116_
  (
    .in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_116_out)
  );


  direct_interc
  direct_interc_117_
  (
    .in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_117_out)
  );


  direct_interc
  direct_interc_118_
  (
    .in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_118_out)
  );


  direct_interc
  direct_interc_119_
  (
    .in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_119_out)
  );


  direct_interc
  direct_interc_120_
  (
    .in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_120_out)
  );


  direct_interc
  direct_interc_121_
  (
    .in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_121_out)
  );


  direct_interc
  direct_interc_122_
  (
    .in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_122_out)
  );


  direct_interc
  direct_interc_123_
  (
    .in(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_123_out)
  );


  direct_interc
  direct_interc_124_
  (
    .in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_124_out)
  );


  direct_interc
  direct_interc_125_
  (
    .in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_125_out)
  );


  direct_interc
  direct_interc_126_
  (
    .in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_126_out)
  );


  direct_interc
  direct_interc_127_
  (
    .in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_127_out)
  );


  direct_interc
  direct_interc_128_
  (
    .in(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_128_out)
  );


  direct_interc
  direct_interc_129_
  (
    .in(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_129_out)
  );


  direct_interc
  direct_interc_130_
  (
    .in(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_130_out)
  );


  direct_interc
  direct_interc_131_
  (
    .in(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_131_out)
  );


  direct_interc
  direct_interc_132_
  (
    .in(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_132_out)
  );


  direct_interc
  direct_interc_133_
  (
    .in(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_133_out)
  );


  direct_interc
  direct_interc_134_
  (
    .in(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_134_out)
  );


  direct_interc
  direct_interc_135_
  (
    .in(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_135_out)
  );


  direct_interc
  direct_interc_136_
  (
    .in(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_136_out)
  );


  direct_interc
  direct_interc_137_
  (
    .in(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_137_out)
  );


  direct_interc
  direct_interc_138_
  (
    .in(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_138_out)
  );


  direct_interc
  direct_interc_139_
  (
    .in(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_139_out)
  );


  direct_interc
  direct_interc_140_
  (
    .in(grid_clb_81_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_140_out)
  );


  direct_interc
  direct_interc_141_
  (
    .in(grid_clb_83_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_141_out)
  );


  direct_interc
  direct_interc_142_
  (
    .in(grid_clb_84_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_142_out)
  );


  direct_interc
  direct_interc_143_
  (
    .in(grid_clb_85_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_143_out)
  );


  direct_interc
  direct_interc_144_
  (
    .in(grid_clb_86_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_144_out)
  );


  direct_interc
  direct_interc_145_
  (
    .in(grid_clb_87_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_145_out)
  );


  direct_interc
  direct_interc_146_
  (
    .in(grid_clb_89_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_146_out)
  );


  direct_interc
  direct_interc_147_
  (
    .in(grid_clb_91_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_147_out)
  );


  direct_interc
  direct_interc_148_
  (
    .in(grid_clb_93_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_148_out)
  );


  direct_interc
  direct_interc_149_
  (
    .in(grid_clb_94_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_149_out)
  );


  direct_interc
  direct_interc_150_
  (
    .in(grid_clb_95_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_150_out)
  );


  direct_interc
  direct_interc_151_
  (
    .in(grid_clb_96_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_151_out)
  );


  direct_interc
  direct_interc_152_
  (
    .in(grid_clb_97_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_152_out)
  );


  direct_interc
  direct_interc_153_
  (
    .in(grid_clb_99_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_153_out)
  );


  direct_interc
  direct_interc_154_
  (
    .in(grid_clb_101_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_154_out)
  );


  direct_interc
  direct_interc_155_
  (
    .in(grid_clb_103_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_155_out)
  );


  direct_interc
  direct_interc_156_
  (
    .in(grid_clb_104_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_156_out)
  );


  direct_interc
  direct_interc_157_
  (
    .in(grid_clb_105_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_157_out)
  );


  direct_interc
  direct_interc_158_
  (
    .in(grid_clb_106_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_158_out)
  );


  direct_interc
  direct_interc_159_
  (
    .in(grid_clb_107_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_159_out)
  );


  direct_interc
  direct_interc_160_
  (
    .in(grid_clb_109_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_160_out)
  );


  direct_interc
  direct_interc_161_
  (
    .in(grid_clb_111_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_161_out)
  );


  direct_interc
  direct_interc_162_
  (
    .in(grid_clb_113_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_162_out)
  );


  direct_interc
  direct_interc_163_
  (
    .in(grid_clb_114_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_163_out)
  );


  direct_interc
  direct_interc_164_
  (
    .in(grid_clb_115_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_164_out)
  );


  direct_interc
  direct_interc_165_
  (
    .in(grid_clb_116_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_165_out)
  );


  direct_interc
  direct_interc_166_
  (
    .in(grid_clb_117_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_166_out)
  );


  direct_interc
  direct_interc_167_
  (
    .in(grid_clb_119_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_167_out)
  );


  direct_interc
  direct_interc_168_
  (
    .in(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_168_out)
  );


  direct_interc
  direct_interc_169_
  (
    .in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_169_out)
  );


  direct_interc
  direct_interc_170_
  (
    .in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_170_out)
  );


  direct_interc
  direct_interc_171_
  (
    .in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_171_out)
  );


  direct_interc
  direct_interc_172_
  (
    .in(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_172_out)
  );


  direct_interc
  direct_interc_173_
  (
    .in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_173_out)
  );


  direct_interc
  direct_interc_174_
  (
    .in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_174_out)
  );


  direct_interc
  direct_interc_175_
  (
    .in(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_175_out)
  );


  direct_interc
  direct_interc_176_
  (
    .in(grid_clb_80_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_176_out)
  );


  direct_interc
  direct_interc_177_
  (
    .in(grid_clb_90_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_177_out)
  );


  direct_interc
  direct_interc_178_
  (
    .in(grid_clb_100_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
    .out(direct_interc_178_out)
  );


endmodule

