

module frac_mult_18_18
(
  input [0:17] A,
  input [0:17] B,
  output [0:35] Y,
  input [0:0] MODE
);

  wire MODE_0_0;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  assign MODE_0_0 = MODE[0];

  sky130_fd_sc_hd__mux2i_1
  U38
  (
    .A0(n24),
    .A1(n25),
    .S(MODE_0_0),
    .Y(Y[9])
  );


  sky130_fd_sc_hd__xnor2_1
  U39
  (
    .A(n26),
    .B(n27),
    .Y(n25)
  );


  sky130_fd_sc_hd__xnor2_1
  U40
  (
    .A(n28),
    .B(n29),
    .Y(n27)
  );


  sky130_fd_sc_hd__xnor2_1
  U41
  (
    .A(n30),
    .B(n31),
    .Y(n24)
  );


  sky130_fd_sc_hd__xor2_1
  U42
  (
    .A(n32),
    .B(n33),
    .X(n31)
  );


  sky130_fd_sc_hd__mux2i_1
  U43
  (
    .A0(n34),
    .A1(n35),
    .S(MODE_0_0),
    .Y(Y[8])
  );


  sky130_fd_sc_hd__xnor2_1
  U44
  (
    .A(n36),
    .B(n37),
    .Y(n35)
  );


  sky130_fd_sc_hd__xor2_1
  U45
  (
    .A(n38),
    .B(n39),
    .X(n37)
  );


  sky130_fd_sc_hd__xnor2_1
  U46
  (
    .A(n40),
    .B(n41),
    .Y(n34)
  );


  sky130_fd_sc_hd__xnor2_1
  U47
  (
    .A(n42),
    .B(n43),
    .Y(n41)
  );


  sky130_fd_sc_hd__mux2i_1
  U48
  (
    .A0(n44),
    .A1(n45),
    .S(MODE_0_0),
    .Y(Y[7])
  );


  sky130_fd_sc_hd__xnor2_1
  U49
  (
    .A(n46),
    .B(n47),
    .Y(n45)
  );


  sky130_fd_sc_hd__xnor2_1
  U50
  (
    .A(n48),
    .B(n49),
    .Y(n46)
  );


  sky130_fd_sc_hd__xnor2_1
  U51
  (
    .A(n50),
    .B(n51),
    .Y(n44)
  );


  sky130_fd_sc_hd__xor2_1
  U52
  (
    .A(n52),
    .B(n53),
    .X(n50)
  );


  sky130_fd_sc_hd__mux2i_1
  U53
  (
    .A0(n54),
    .A1(n55),
    .S(MODE_0_0),
    .Y(Y[6])
  );


  sky130_fd_sc_hd__xnor2_1
  U54
  (
    .A(n56),
    .B(n57),
    .Y(n55)
  );


  sky130_fd_sc_hd__xor2_1
  U55
  (
    .A(n58),
    .B(n59),
    .X(n56)
  );


  sky130_fd_sc_hd__xnor2_1
  U56
  (
    .A(n60),
    .B(n61),
    .Y(n54)
  );


  sky130_fd_sc_hd__xor2_1
  U57
  (
    .A(n62),
    .B(n63),
    .X(n61)
  );


  sky130_fd_sc_hd__mux2i_1
  U58
  (
    .A0(n64),
    .A1(n65),
    .S(MODE_0_0),
    .Y(Y[5])
  );


  sky130_fd_sc_hd__xnor2_1
  U59
  (
    .A(n66),
    .B(n67),
    .Y(n65)
  );


  sky130_fd_sc_hd__xnor2_1
  U60
  (
    .A(n68),
    .B(n69),
    .Y(n67)
  );


  sky130_fd_sc_hd__xnor2_1
  U61
  (
    .A(n70),
    .B(n71),
    .Y(n64)
  );


  sky130_fd_sc_hd__xnor2_1
  U62
  (
    .A(n72),
    .B(n73),
    .Y(n71)
  );


  sky130_fd_sc_hd__mux2i_1
  U63
  (
    .A0(n74),
    .A1(n75),
    .S(MODE_0_0),
    .Y(Y[4])
  );


  sky130_fd_sc_hd__xnor2_1
  U64
  (
    .A(n76),
    .B(n77),
    .Y(n75)
  );


  sky130_fd_sc_hd__xor2_1
  U65
  (
    .A(n78),
    .B(n79),
    .X(n76)
  );


  sky130_fd_sc_hd__xnor2_1
  U66
  (
    .A(n80),
    .B(n81),
    .Y(n74)
  );


  sky130_fd_sc_hd__xor2_1
  U67
  (
    .A(n82),
    .B(n83),
    .X(n80)
  );


  sky130_fd_sc_hd__mux2i_1
  U68
  (
    .A0(n84),
    .A1(n85),
    .S(MODE_0_0),
    .Y(Y[3])
  );


  sky130_fd_sc_hd__xnor2_1
  U69
  (
    .A(n86),
    .B(n87),
    .Y(n85)
  );


  sky130_fd_sc_hd__xor2_1
  U70
  (
    .A(n88),
    .B(n89),
    .X(n87)
  );


  sky130_fd_sc_hd__xnor2_1
  U71
  (
    .A(n90),
    .B(n91),
    .Y(n84)
  );


  sky130_fd_sc_hd__xor2_1
  U72
  (
    .A(n92),
    .B(n93),
    .X(n91)
  );


  sky130_fd_sc_hd__xor2_1
  U73
  (
    .A(A[15]),
    .B(n94),
    .X(Y[35])
  );


  sky130_fd_sc_hd__xor2_1
  U74
  (
    .A(n95),
    .B(n96),
    .X(Y[34])
  );


  sky130_fd_sc_hd__nor2b_1
  U75
  (
    .B_N(n94),
    .A(n97),
    .Y(n96)
  );


  sky130_fd_sc_hd__xor2_1
  U76
  (
    .A(n98),
    .B(n99),
    .X(Y[33])
  );


  sky130_fd_sc_hd__xnor2_1
  U77
  (
    .A(n100),
    .B(n101),
    .Y(Y[32])
  );


  sky130_fd_sc_hd__nor2_1
  U78
  (
    .A(n102),
    .B(n103),
    .Y(n100)
  );


  sky130_fd_sc_hd__xor2_1
  U79
  (
    .A(n104),
    .B(n105),
    .X(Y[31])
  );


  sky130_fd_sc_hd__xnor2_1
  U80
  (
    .A(n106),
    .B(n107),
    .Y(n104)
  );


  sky130_fd_sc_hd__xor2_1
  U81
  (
    .A(n108),
    .B(n109),
    .X(Y[30])
  );


  sky130_fd_sc_hd__xnor2_1
  U82
  (
    .A(n110),
    .B(n111),
    .Y(n108)
  );


  sky130_fd_sc_hd__mux2i_1
  U83
  (
    .A0(n112),
    .A1(n113),
    .S(MODE_0_0),
    .Y(Y[2])
  );


  sky130_fd_sc_hd__xnor2_1
  U84
  (
    .A(n114),
    .B(n115),
    .Y(n113)
  );


  sky130_fd_sc_hd__xor2_1
  U85
  (
    .A(n116),
    .B(n117),
    .X(n114)
  );


  sky130_fd_sc_hd__xnor2_1
  U86
  (
    .A(n118),
    .B(n119),
    .Y(n112)
  );


  sky130_fd_sc_hd__xnor2_1
  U87
  (
    .A(n120),
    .B(n121),
    .Y(n119)
  );


  sky130_fd_sc_hd__xor2_1
  U88
  (
    .A(n122),
    .B(n123),
    .X(Y[29])
  );


  sky130_fd_sc_hd__xnor2_1
  U89
  (
    .A(n124),
    .B(n125),
    .Y(n122)
  );


  sky130_fd_sc_hd__xor2_1
  U90
  (
    .A(n126),
    .B(n127),
    .X(Y[28])
  );


  sky130_fd_sc_hd__xnor2_1
  U91
  (
    .A(n128),
    .B(n129),
    .Y(n126)
  );


  sky130_fd_sc_hd__xor2_1
  U92
  (
    .A(n130),
    .B(n131),
    .X(Y[27])
  );


  sky130_fd_sc_hd__xnor2_1
  U93
  (
    .A(n132),
    .B(n133),
    .Y(n130)
  );


  sky130_fd_sc_hd__xor2_1
  U94
  (
    .A(n134),
    .B(n135),
    .X(Y[26])
  );


  sky130_fd_sc_hd__xnor2_1
  U95
  (
    .A(n136),
    .B(n137),
    .Y(n134)
  );


  sky130_fd_sc_hd__xor2_1
  U96
  (
    .A(n138),
    .B(n139),
    .X(Y[25])
  );


  sky130_fd_sc_hd__xnor2_1
  U97
  (
    .A(n140),
    .B(n141),
    .Y(n138)
  );


  sky130_fd_sc_hd__xor2_1
  U98
  (
    .A(n142),
    .B(n143),
    .X(Y[24])
  );


  sky130_fd_sc_hd__xnor2_1
  U99
  (
    .A(n144),
    .B(n145),
    .Y(n142)
  );


  sky130_fd_sc_hd__xor2_1
  U100
  (
    .A(n146),
    .B(n147),
    .X(Y[23])
  );


  sky130_fd_sc_hd__xnor2_1
  U101
  (
    .A(n148),
    .B(n149),
    .Y(n146)
  );


  sky130_fd_sc_hd__xor2_1
  U102
  (
    .A(n150),
    .B(n151),
    .X(Y[22])
  );


  sky130_fd_sc_hd__xnor2_1
  U103
  (
    .A(n152),
    .B(n153),
    .Y(n150)
  );


  sky130_fd_sc_hd__xor2_1
  U104
  (
    .A(n154),
    .B(n155),
    .X(Y[21])
  );


  sky130_fd_sc_hd__xnor2_1
  U105
  (
    .A(n156),
    .B(n157),
    .Y(n154)
  );


  sky130_fd_sc_hd__xor2_1
  U106
  (
    .A(n158),
    .B(n159),
    .X(Y[20])
  );


  sky130_fd_sc_hd__xnor2_1
  U107
  (
    .A(n160),
    .B(n161),
    .Y(n158)
  );


  sky130_fd_sc_hd__mux2i_1
  U108
  (
    .A0(n162),
    .A1(n163),
    .S(MODE_0_0),
    .Y(Y[1])
  );


  sky130_fd_sc_hd__xnor2_1
  U109
  (
    .A(n164),
    .B(n165),
    .Y(n163)
  );


  sky130_fd_sc_hd__xor2_1
  U110
  (
    .A(n166),
    .B(n167),
    .X(n165)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U111
  (
    .B1(n168),
    .B2(n169),
    .A1_N(n170),
    .A2_N(n171),
    .Y(n167)
  );


  sky130_fd_sc_hd__nor2_1
  U112
  (
    .A(n168),
    .B(n169),
    .Y(n170)
  );


  sky130_fd_sc_hd__o22ai_1
  U113
  (
    .A1(n117),
    .A2(n172),
    .B1(n173),
    .B2(n115),
    .Y(n166)
  );


  sky130_fd_sc_hd__and2_0
  U114
  (
    .A(n117),
    .B(n172),
    .X(n173)
  );


  sky130_fd_sc_hd__clkinv_1
  U115
  (
    .A(n116),
    .Y(n172)
  );


  sky130_fd_sc_hd__o22ai_1
  U116
  (
    .A1(n89),
    .A2(n174),
    .B1(n175),
    .B2(n86),
    .Y(n116)
  );


  sky130_fd_sc_hd__and2_0
  U117
  (
    .A(n89),
    .B(n174),
    .X(n175)
  );


  sky130_fd_sc_hd__clkinv_1
  U118
  (
    .A(n88),
    .Y(n174)
  );


  sky130_fd_sc_hd__o22ai_1
  U119
  (
    .A1(n79),
    .A2(n176),
    .B1(n177),
    .B2(n77),
    .Y(n88)
  );


  sky130_fd_sc_hd__nor2_1
  U120
  (
    .A(n178),
    .B(n78),
    .Y(n177)
  );


  sky130_fd_sc_hd__clkinv_1
  U121
  (
    .A(n176),
    .Y(n78)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U122
  (
    .B1(n69),
    .B2(n68),
    .A1_N(n179),
    .A2_N(n66),
    .Y(n176)
  );


  sky130_fd_sc_hd__nor2_1
  U123
  (
    .A(n69),
    .B(n68),
    .Y(n179)
  );


  sky130_fd_sc_hd__o22ai_1
  U124
  (
    .A1(n59),
    .A2(n180),
    .B1(n181),
    .B2(n57),
    .Y(n68)
  );


  sky130_fd_sc_hd__nor2_1
  U125
  (
    .A(n182),
    .B(n58),
    .Y(n181)
  );


  sky130_fd_sc_hd__clkinv_1
  U126
  (
    .A(n180),
    .Y(n58)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U127
  (
    .B1(n49),
    .B2(n48),
    .A1_N(n183),
    .A2_N(n47),
    .Y(n180)
  );


  sky130_fd_sc_hd__nor2_1
  U128
  (
    .A(n49),
    .B(n48),
    .Y(n183)
  );


  sky130_fd_sc_hd__o22ai_1
  U129
  (
    .A1(n39),
    .A2(n184),
    .B1(n185),
    .B2(n36),
    .Y(n48)
  );


  sky130_fd_sc_hd__nor2_1
  U130
  (
    .A(n186),
    .B(n38),
    .Y(n185)
  );


  sky130_fd_sc_hd__clkinv_1
  U131
  (
    .A(n184),
    .Y(n38)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U132
  (
    .B1(n29),
    .B2(n28),
    .A1_N(n187),
    .A2_N(n26),
    .Y(n184)
  );


  sky130_fd_sc_hd__nor2_1
  U133
  (
    .A(n29),
    .B(n28),
    .Y(n187)
  );


  sky130_fd_sc_hd__o22ai_1
  U134
  (
    .A1(n188),
    .A2(n189),
    .B1(n190),
    .B2(n191),
    .Y(n28)
  );


  sky130_fd_sc_hd__nor2_1
  U135
  (
    .A(n192),
    .B(n193),
    .Y(n190)
  );


  sky130_fd_sc_hd__clkinv_1
  U136
  (
    .A(n192),
    .Y(n189)
  );


  sky130_fd_sc_hd__o22ai_1
  U137
  (
    .A1(n194),
    .A2(n195),
    .B1(n196),
    .B2(n197),
    .Y(n29)
  );


  sky130_fd_sc_hd__nor2_1
  U138
  (
    .A(n198),
    .B(n199),
    .Y(n196)
  );


  sky130_fd_sc_hd__clkinv_1
  U139
  (
    .A(n186),
    .Y(n39)
  );


  sky130_fd_sc_hd__o22ai_1
  U140
  (
    .A1(n200),
    .A2(n201),
    .B1(n202),
    .B2(n203),
    .Y(n186)
  );


  sky130_fd_sc_hd__nor2_1
  U141
  (
    .A(n204),
    .B(n205),
    .Y(n202)
  );


  sky130_fd_sc_hd__o22ai_1
  U142
  (
    .A1(n206),
    .A2(n207),
    .B1(n208),
    .B2(n209),
    .Y(n49)
  );


  sky130_fd_sc_hd__and2_0
  U143
  (
    .A(n207),
    .B(n206),
    .X(n208)
  );


  sky130_fd_sc_hd__clkinv_1
  U144
  (
    .A(n182),
    .Y(n59)
  );


  sky130_fd_sc_hd__o22ai_1
  U145
  (
    .A1(n210),
    .A2(n211),
    .B1(n212),
    .B2(n213),
    .Y(n182)
  );


  sky130_fd_sc_hd__and2_0
  U146
  (
    .A(n211),
    .B(n210),
    .X(n212)
  );


  sky130_fd_sc_hd__o22ai_1
  U147
  (
    .A1(n214),
    .A2(n215),
    .B1(n216),
    .B2(n217),
    .Y(n69)
  );


  sky130_fd_sc_hd__and2_0
  U148
  (
    .A(n215),
    .B(n214),
    .X(n216)
  );


  sky130_fd_sc_hd__clkinv_1
  U149
  (
    .A(n178),
    .Y(n79)
  );


  sky130_fd_sc_hd__o22ai_1
  U150
  (
    .A1(n218),
    .A2(n219),
    .B1(n220),
    .B2(n221),
    .Y(n178)
  );


  sky130_fd_sc_hd__and2_0
  U151
  (
    .A(n219),
    .B(n218),
    .X(n220)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U152
  (
    .B1(n222),
    .B2(n223),
    .A1_N(n224),
    .A2_N(n225),
    .Y(n89)
  );


  sky130_fd_sc_hd__nor2_1
  U153
  (
    .A(n222),
    .B(n223),
    .Y(n224)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U154
  (
    .B1(n226),
    .B2(n227),
    .A1_N(n228),
    .A2_N(n229),
    .Y(n117)
  );


  sky130_fd_sc_hd__nor2_1
  U155
  (
    .A(n226),
    .B(n227),
    .Y(n228)
  );


  sky130_fd_sc_hd__xnor2_1
  U156
  (
    .A(n230),
    .B(n231),
    .Y(n162)
  );


  sky130_fd_sc_hd__xor2_1
  U157
  (
    .A(n232),
    .B(n233),
    .X(n230)
  );


  sky130_fd_sc_hd__o22a_1
  U158
  (
    .A1(n234),
    .A2(n235),
    .B1(n236),
    .B2(n237),
    .X(n233)
  );


  sky130_fd_sc_hd__nor2b_1
  U159
  (
    .B_N(n235),
    .A(n238),
    .Y(n237)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U160
  (
    .B1(n239),
    .B2(n118),
    .A1_N(n121),
    .A2_N(n120),
    .Y(n232)
  );


  sky130_fd_sc_hd__nor2_1
  U161
  (
    .A(n121),
    .B(n120),
    .Y(n239)
  );


  sky130_fd_sc_hd__o22ai_1
  U162
  (
    .A1(n93),
    .A2(n240),
    .B1(n241),
    .B2(n90),
    .Y(n120)
  );


  sky130_fd_sc_hd__and2_0
  U163
  (
    .A(n93),
    .B(n240),
    .X(n241)
  );


  sky130_fd_sc_hd__clkinv_1
  U164
  (
    .A(n92),
    .Y(n240)
  );


  sky130_fd_sc_hd__o22ai_1
  U165
  (
    .A1(n83),
    .A2(n242),
    .B1(n243),
    .B2(n81),
    .Y(n92)
  );


  sky130_fd_sc_hd__nor2_1
  U166
  (
    .A(n244),
    .B(n82),
    .Y(n243)
  );


  sky130_fd_sc_hd__clkinv_1
  U167
  (
    .A(n242),
    .Y(n82)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U168
  (
    .B1(n73),
    .B2(n72),
    .A1_N(n245),
    .A2_N(n70),
    .Y(n242)
  );


  sky130_fd_sc_hd__nor2_1
  U169
  (
    .A(n73),
    .B(n72),
    .Y(n245)
  );


  sky130_fd_sc_hd__o22ai_1
  U170
  (
    .A1(n63),
    .A2(n246),
    .B1(n247),
    .B2(n60),
    .Y(n72)
  );


  sky130_fd_sc_hd__and2_0
  U171
  (
    .A(n63),
    .B(n246),
    .X(n247)
  );


  sky130_fd_sc_hd__clkinv_1
  U172
  (
    .A(n62),
    .Y(n246)
  );


  sky130_fd_sc_hd__o22ai_1
  U173
  (
    .A1(n53),
    .A2(n248),
    .B1(n249),
    .B2(n51),
    .Y(n62)
  );


  sky130_fd_sc_hd__nor2_1
  U174
  (
    .A(n250),
    .B(n52),
    .Y(n249)
  );


  sky130_fd_sc_hd__clkinv_1
  U175
  (
    .A(n248),
    .Y(n52)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U176
  (
    .B1(n43),
    .B2(n42),
    .A1_N(n251),
    .A2_N(n40),
    .Y(n248)
  );


  sky130_fd_sc_hd__nor2_1
  U177
  (
    .A(n43),
    .B(n42),
    .Y(n251)
  );


  sky130_fd_sc_hd__o22ai_1
  U178
  (
    .A1(n33),
    .A2(n252),
    .B1(n253),
    .B2(n30),
    .Y(n42)
  );


  sky130_fd_sc_hd__and2_0
  U179
  (
    .A(n33),
    .B(n252),
    .X(n253)
  );


  sky130_fd_sc_hd__clkinv_1
  U180
  (
    .A(n32),
    .Y(n252)
  );


  sky130_fd_sc_hd__o22ai_1
  U181
  (
    .A1(n254),
    .A2(n255),
    .B1(n256),
    .B2(n257),
    .Y(n32)
  );


  sky130_fd_sc_hd__nor2_1
  U182
  (
    .A(n258),
    .B(n259),
    .Y(n256)
  );


  sky130_fd_sc_hd__clkinv_1
  U183
  (
    .A(n258),
    .Y(n255)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U184
  (
    .B1(n260),
    .B2(n261),
    .A1_N(n262),
    .A2_N(n263),
    .Y(n33)
  );


  sky130_fd_sc_hd__nor2_1
  U185
  (
    .A(n261),
    .B(n260),
    .Y(n262)
  );


  sky130_fd_sc_hd__o22ai_1
  U186
  (
    .A1(n264),
    .A2(n265),
    .B1(n266),
    .B2(n267),
    .Y(n43)
  );


  sky130_fd_sc_hd__and2_0
  U187
  (
    .A(n265),
    .B(n264),
    .X(n266)
  );


  sky130_fd_sc_hd__clkinv_1
  U188
  (
    .A(n250),
    .Y(n53)
  );


  sky130_fd_sc_hd__o22ai_1
  U189
  (
    .A1(n268),
    .A2(n269),
    .B1(n270),
    .B2(n271),
    .Y(n250)
  );


  sky130_fd_sc_hd__and2_0
  U190
  (
    .A(n269),
    .B(n268),
    .X(n270)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U191
  (
    .B1(n272),
    .B2(n273),
    .A1_N(n274),
    .A2_N(n275),
    .Y(n63)
  );


  sky130_fd_sc_hd__nor2_1
  U192
  (
    .A(n273),
    .B(n272),
    .Y(n274)
  );


  sky130_fd_sc_hd__o22ai_1
  U193
  (
    .A1(n276),
    .A2(n277),
    .B1(n278),
    .B2(n279),
    .Y(n73)
  );


  sky130_fd_sc_hd__and2_0
  U194
  (
    .A(n277),
    .B(n276),
    .X(n278)
  );


  sky130_fd_sc_hd__clkinv_1
  U195
  (
    .A(n244),
    .Y(n83)
  );


  sky130_fd_sc_hd__o22ai_1
  U196
  (
    .A1(n280),
    .A2(n281),
    .B1(n282),
    .B2(n283),
    .Y(n244)
  );


  sky130_fd_sc_hd__and2_0
  U197
  (
    .A(n281),
    .B(n280),
    .X(n282)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U198
  (
    .B1(n284),
    .B2(n285),
    .A1_N(n286),
    .A2_N(n287),
    .Y(n93)
  );


  sky130_fd_sc_hd__nor2_1
  U199
  (
    .A(n285),
    .B(n284),
    .Y(n286)
  );


  sky130_fd_sc_hd__o22ai_1
  U200
  (
    .A1(n288),
    .A2(n289),
    .B1(n290),
    .B2(n291),
    .Y(n121)
  );


  sky130_fd_sc_hd__and2_0
  U201
  (
    .A(n289),
    .B(n288),
    .X(n290)
  );


  sky130_fd_sc_hd__xor2_1
  U202
  (
    .A(n292),
    .B(n293),
    .X(Y[19])
  );


  sky130_fd_sc_hd__xnor2_1
  U203
  (
    .A(n294),
    .B(n295),
    .Y(n292)
  );


  sky130_fd_sc_hd__xor2_1
  U204
  (
    .A(n296),
    .B(n297),
    .X(Y[18])
  );


  sky130_fd_sc_hd__xnor2_1
  U205
  (
    .A(n298),
    .B(n299),
    .Y(n296)
  );


  sky130_fd_sc_hd__o31ai_1
  U206
  (
    .A1(n300),
    .A2(n301),
    .A3(n302),
    .B1(n303),
    .Y(Y[17])
  );


  sky130_fd_sc_hd__xor2_1
  U207
  (
    .A(n304),
    .B(n305),
    .X(n303)
  );


  sky130_fd_sc_hd__xor2_1
  U208
  (
    .A(n306),
    .B(n307),
    .X(n305)
  );


  sky130_fd_sc_hd__o21ai_0
  U209
  (
    .A1(n308),
    .A2(n300),
    .B1(n309),
    .Y(Y[16])
  );


  sky130_fd_sc_hd__xnor2_1
  U210
  (
    .A(n310),
    .B(n311),
    .Y(n309)
  );


  sky130_fd_sc_hd__xnor2_1
  U211
  (
    .A(n312),
    .B(n313),
    .Y(n310)
  );


  sky130_fd_sc_hd__xor2_1
  U212
  (
    .A(n314),
    .B(n315),
    .X(n308)
  );


  sky130_fd_sc_hd__o21ai_0
  U213
  (
    .A1(n300),
    .A2(n316),
    .B1(n317),
    .Y(Y[15])
  );


  sky130_fd_sc_hd__xnor2_1
  U214
  (
    .A(n318),
    .B(n319),
    .Y(n317)
  );


  sky130_fd_sc_hd__xnor2_1
  U215
  (
    .A(n320),
    .B(n321),
    .Y(n319)
  );


  sky130_fd_sc_hd__xor2_1
  U216
  (
    .A(n322),
    .B(n323),
    .X(n316)
  );


  sky130_fd_sc_hd__nand2_1
  U217
  (
    .A(n324),
    .B(n325),
    .Y(n322)
  );


  sky130_fd_sc_hd__o21ai_0
  U218
  (
    .A1(n300),
    .A2(n326),
    .B1(n327),
    .Y(Y[14])
  );


  sky130_fd_sc_hd__xnor2_1
  U219
  (
    .A(n328),
    .B(n329),
    .Y(n327)
  );


  sky130_fd_sc_hd__xor2_1
  U220
  (
    .A(n330),
    .B(n331),
    .X(n329)
  );


  sky130_fd_sc_hd__xor2_1
  U221
  (
    .A(n332),
    .B(n333),
    .X(n326)
  );


  sky130_fd_sc_hd__xor2_1
  U222
  (
    .A(n334),
    .B(n335),
    .X(n333)
  );


  sky130_fd_sc_hd__o21ai_0
  U223
  (
    .A1(n300),
    .A2(n336),
    .B1(n337),
    .Y(Y[13])
  );


  sky130_fd_sc_hd__xnor2_1
  U224
  (
    .A(n338),
    .B(n339),
    .Y(n337)
  );


  sky130_fd_sc_hd__xnor2_1
  U225
  (
    .A(n340),
    .B(n341),
    .Y(n339)
  );


  sky130_fd_sc_hd__xor2_1
  U226
  (
    .A(n342),
    .B(n343),
    .X(n336)
  );


  sky130_fd_sc_hd__xor2_1
  U227
  (
    .A(n344),
    .B(n345),
    .X(n343)
  );


  sky130_fd_sc_hd__o21ai_0
  U228
  (
    .A1(n300),
    .A2(n346),
    .B1(n347),
    .Y(Y[12])
  );


  sky130_fd_sc_hd__xnor2_1
  U229
  (
    .A(n348),
    .B(n349),
    .Y(n347)
  );


  sky130_fd_sc_hd__xor2_1
  U230
  (
    .A(n350),
    .B(n351),
    .X(n348)
  );


  sky130_fd_sc_hd__xor2_1
  U231
  (
    .A(n352),
    .B(n353),
    .X(n346)
  );


  sky130_fd_sc_hd__xor2_1
  U232
  (
    .A(n354),
    .B(n355),
    .X(n353)
  );


  sky130_fd_sc_hd__mux2i_1
  U233
  (
    .A0(n356),
    .A1(n357),
    .S(MODE_0_0),
    .Y(Y[11])
  );


  sky130_fd_sc_hd__xnor2_1
  U234
  (
    .A(n358),
    .B(n359),
    .Y(n357)
  );


  sky130_fd_sc_hd__xnor2_1
  U235
  (
    .A(n360),
    .B(n361),
    .Y(n359)
  );


  sky130_fd_sc_hd__xnor2_1
  U236
  (
    .A(n362),
    .B(n363),
    .Y(n356)
  );


  sky130_fd_sc_hd__xnor2_1
  U237
  (
    .A(n364),
    .B(n365),
    .Y(n363)
  );


  sky130_fd_sc_hd__mux2i_1
  U238
  (
    .A0(n366),
    .A1(n367),
    .S(MODE_0_0),
    .Y(Y[10])
  );


  sky130_fd_sc_hd__xnor2_1
  U239
  (
    .A(n191),
    .B(n368),
    .Y(n367)
  );


  sky130_fd_sc_hd__xor2_1
  U240
  (
    .A(n192),
    .B(n188),
    .X(n368)
  );


  sky130_fd_sc_hd__clkinv_1
  U241
  (
    .A(n193),
    .Y(n188)
  );


  sky130_fd_sc_hd__o22ai_1
  U242
  (
    .A1(n369),
    .A2(n370),
    .B1(n371),
    .B2(n372),
    .Y(n193)
  );


  sky130_fd_sc_hd__nor2_1
  U243
  (
    .A(n373),
    .B(n374),
    .Y(n371)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U244
  (
    .B1(n375),
    .B2(n358),
    .A1_N(n361),
    .A2_N(n360),
    .Y(n192)
  );


  sky130_fd_sc_hd__nor2_1
  U245
  (
    .A(n360),
    .B(n361),
    .Y(n375)
  );


  sky130_fd_sc_hd__o22ai_1
  U246
  (
    .A1(n376),
    .A2(n377),
    .B1(n378),
    .B2(n379),
    .Y(n361)
  );


  sky130_fd_sc_hd__nor2_1
  U247
  (
    .A(n380),
    .B(n381),
    .Y(n378)
  );


  sky130_fd_sc_hd__o22ai_1
  U248
  (
    .A1(n354),
    .A2(n355),
    .B1(n382),
    .B2(n352),
    .Y(n360)
  );


  sky130_fd_sc_hd__nor2b_1
  U249
  (
    .B_N(n354),
    .A(n383),
    .Y(n382)
  );


  sky130_fd_sc_hd__clkinv_1
  U250
  (
    .A(n383),
    .Y(n355)
  );


  sky130_fd_sc_hd__o22ai_1
  U251
  (
    .A1(n384),
    .A2(n385),
    .B1(n386),
    .B2(n342),
    .Y(n383)
  );


  sky130_fd_sc_hd__nor2_1
  U252
  (
    .A(n345),
    .B(n344),
    .Y(n386)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U253
  (
    .B1(n387),
    .B2(n388),
    .A1_N(n389),
    .A2_N(n390),
    .Y(n354)
  );


  sky130_fd_sc_hd__nor2_1
  U254
  (
    .A(n388),
    .B(n387),
    .Y(n389)
  );


  sky130_fd_sc_hd__xnor2_1
  U255
  (
    .A(n391),
    .B(n257),
    .Y(n366)
  );


  sky130_fd_sc_hd__xor2_1
  U256
  (
    .A(n258),
    .B(n254),
    .X(n391)
  );


  sky130_fd_sc_hd__clkinv_1
  U257
  (
    .A(n259),
    .Y(n254)
  );


  sky130_fd_sc_hd__o22ai_1
  U258
  (
    .A1(n392),
    .A2(n393),
    .B1(n394),
    .B2(n395),
    .Y(n259)
  );


  sky130_fd_sc_hd__nor2_1
  U259
  (
    .A(n396),
    .B(n397),
    .Y(n394)
  );


  sky130_fd_sc_hd__clkinv_1
  U260
  (
    .A(n396),
    .Y(n393)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U261
  (
    .B1(n398),
    .B2(n362),
    .A1_N(n365),
    .A2_N(n364),
    .Y(n258)
  );


  sky130_fd_sc_hd__nor2_1
  U262
  (
    .A(n364),
    .B(n365),
    .Y(n398)
  );


  sky130_fd_sc_hd__o22ai_1
  U263
  (
    .A1(n399),
    .A2(n400),
    .B1(n401),
    .B2(n402),
    .Y(n365)
  );


  sky130_fd_sc_hd__and2_0
  U264
  (
    .A(n400),
    .B(n399),
    .X(n401)
  );


  sky130_fd_sc_hd__o22ai_1
  U265
  (
    .A1(n351),
    .A2(n403),
    .B1(n404),
    .B2(n349),
    .Y(n364)
  );


  sky130_fd_sc_hd__nor2_1
  U266
  (
    .A(n350),
    .B(n405),
    .Y(n404)
  );


  sky130_fd_sc_hd__clkinv_1
  U267
  (
    .A(n350),
    .Y(n403)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U268
  (
    .B1(n406),
    .B2(n338),
    .A1_N(n341),
    .A2_N(n340),
    .Y(n350)
  );


  sky130_fd_sc_hd__nor2_1
  U269
  (
    .A(n340),
    .B(n341),
    .Y(n406)
  );


  sky130_fd_sc_hd__o22ai_1
  U270
  (
    .A1(n407),
    .A2(n408),
    .B1(n409),
    .B2(n410),
    .Y(n341)
  );


  sky130_fd_sc_hd__and2_0
  U271
  (
    .A(n408),
    .B(n407),
    .X(n409)
  );


  sky130_fd_sc_hd__o22ai_1
  U272
  (
    .A1(n331),
    .A2(n411),
    .B1(n412),
    .B2(n328),
    .Y(n340)
  );


  sky130_fd_sc_hd__nor2_1
  U273
  (
    .A(n330),
    .B(n413),
    .Y(n412)
  );


  sky130_fd_sc_hd__clkinv_1
  U274
  (
    .A(n330),
    .Y(n411)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U275
  (
    .B1(n414),
    .B2(n318),
    .A1_N(n321),
    .A2_N(n320),
    .Y(n330)
  );


  sky130_fd_sc_hd__nor2_1
  U276
  (
    .A(n320),
    .B(n321),
    .Y(n414)
  );


  sky130_fd_sc_hd__o22ai_1
  U277
  (
    .A1(n415),
    .A2(n416),
    .B1(n417),
    .B2(n418),
    .Y(n321)
  );


  sky130_fd_sc_hd__and2_0
  U278
  (
    .A(n416),
    .B(n415),
    .X(n417)
  );


  sky130_fd_sc_hd__o22ai_1
  U279
  (
    .A1(n312),
    .A2(n313),
    .B1(n419),
    .B2(n311),
    .Y(n320)
  );


  sky130_fd_sc_hd__and2_0
  U280
  (
    .A(n313),
    .B(n312),
    .X(n419)
  );


  sky130_fd_sc_hd__xnor2_1
  U281
  (
    .A(n420),
    .B(A[15]),
    .Y(n313)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U282
  (
    .B1(n306),
    .B2(n307),
    .A1_N(n421),
    .A2_N(n304),
    .Y(n312)
  );


  sky130_fd_sc_hd__nor2_1
  U283
  (
    .A(n307),
    .B(n306),
    .Y(n421)
  );


  sky130_fd_sc_hd__xor2_1
  U284
  (
    .A(n97),
    .B(n422),
    .X(n307)
  );


  sky130_fd_sc_hd__o22ai_1
  U285
  (
    .A1(n298),
    .A2(n299),
    .B1(n423),
    .B2(n297),
    .Y(n306)
  );


  sky130_fd_sc_hd__and2_0
  U286
  (
    .A(n299),
    .B(n298),
    .X(n423)
  );


  sky130_fd_sc_hd__xnor2_1
  U287
  (
    .A(n97),
    .B(n424),
    .Y(n299)
  );


  sky130_fd_sc_hd__o22a_1
  U288
  (
    .A1(n294),
    .A2(n295),
    .B1(n425),
    .B2(n293),
    .X(n298)
  );


  sky130_fd_sc_hd__and2_0
  U289
  (
    .A(n295),
    .B(n294),
    .X(n425)
  );


  sky130_fd_sc_hd__xnor2_1
  U290
  (
    .A(n97),
    .B(n426),
    .Y(n295)
  );


  sky130_fd_sc_hd__o22a_1
  U291
  (
    .A1(n160),
    .A2(n161),
    .B1(n427),
    .B2(n159),
    .X(n294)
  );


  sky130_fd_sc_hd__and2_0
  U292
  (
    .A(n161),
    .B(n160),
    .X(n427)
  );


  sky130_fd_sc_hd__xnor2_1
  U293
  (
    .A(n97),
    .B(n428),
    .Y(n161)
  );


  sky130_fd_sc_hd__o22a_1
  U294
  (
    .A1(n156),
    .A2(n157),
    .B1(n429),
    .B2(n155),
    .X(n160)
  );


  sky130_fd_sc_hd__and2_0
  U295
  (
    .A(n157),
    .B(n156),
    .X(n429)
  );


  sky130_fd_sc_hd__xnor2_1
  U296
  (
    .A(n97),
    .B(n430),
    .Y(n157)
  );


  sky130_fd_sc_hd__o22a_1
  U297
  (
    .A1(n152),
    .A2(n153),
    .B1(n431),
    .B2(n151),
    .X(n156)
  );


  sky130_fd_sc_hd__and2_0
  U298
  (
    .A(n153),
    .B(n152),
    .X(n431)
  );


  sky130_fd_sc_hd__xnor2_1
  U299
  (
    .A(n97),
    .B(n432),
    .Y(n153)
  );


  sky130_fd_sc_hd__o22a_1
  U300
  (
    .A1(n148),
    .A2(n149),
    .B1(n433),
    .B2(n147),
    .X(n152)
  );


  sky130_fd_sc_hd__and2_0
  U301
  (
    .A(n149),
    .B(n148),
    .X(n433)
  );


  sky130_fd_sc_hd__xnor2_1
  U302
  (
    .A(n97),
    .B(n434),
    .Y(n149)
  );


  sky130_fd_sc_hd__o22a_1
  U303
  (
    .A1(n144),
    .A2(n145),
    .B1(n435),
    .B2(n143),
    .X(n148)
  );


  sky130_fd_sc_hd__and2_0
  U304
  (
    .A(n145),
    .B(n144),
    .X(n435)
  );


  sky130_fd_sc_hd__xnor2_1
  U305
  (
    .A(n97),
    .B(n436),
    .Y(n145)
  );


  sky130_fd_sc_hd__o22a_1
  U306
  (
    .A1(n140),
    .A2(n141),
    .B1(n437),
    .B2(n139),
    .X(n144)
  );


  sky130_fd_sc_hd__and2_0
  U307
  (
    .A(n141),
    .B(n140),
    .X(n437)
  );


  sky130_fd_sc_hd__xnor2_1
  U308
  (
    .A(n97),
    .B(n438),
    .Y(n141)
  );


  sky130_fd_sc_hd__o22a_1
  U309
  (
    .A1(n136),
    .A2(n137),
    .B1(n439),
    .B2(n135),
    .X(n140)
  );


  sky130_fd_sc_hd__and2_0
  U310
  (
    .A(n137),
    .B(n136),
    .X(n439)
  );


  sky130_fd_sc_hd__xnor2_1
  U311
  (
    .A(n97),
    .B(n440),
    .Y(n137)
  );


  sky130_fd_sc_hd__o22a_1
  U312
  (
    .A1(n132),
    .A2(n133),
    .B1(n441),
    .B2(n131),
    .X(n136)
  );


  sky130_fd_sc_hd__and2_0
  U313
  (
    .A(n133),
    .B(n132),
    .X(n441)
  );


  sky130_fd_sc_hd__xnor2_1
  U314
  (
    .A(n97),
    .B(n442),
    .Y(n133)
  );


  sky130_fd_sc_hd__o22a_1
  U315
  (
    .A1(n128),
    .A2(n129),
    .B1(n443),
    .B2(n127),
    .X(n132)
  );


  sky130_fd_sc_hd__and2_0
  U316
  (
    .A(n129),
    .B(n128),
    .X(n443)
  );


  sky130_fd_sc_hd__xnor2_1
  U317
  (
    .A(n97),
    .B(n444),
    .Y(n129)
  );


  sky130_fd_sc_hd__o22a_1
  U318
  (
    .A1(n124),
    .A2(n125),
    .B1(n445),
    .B2(n123),
    .X(n128)
  );


  sky130_fd_sc_hd__and2_0
  U319
  (
    .A(n125),
    .B(n124),
    .X(n445)
  );


  sky130_fd_sc_hd__xnor2_1
  U320
  (
    .A(n97),
    .B(n446),
    .Y(n125)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U321
  (
    .B1(n111),
    .B2(n110),
    .A1_N(n447),
    .A2_N(n109),
    .Y(n124)
  );


  sky130_fd_sc_hd__nor2_1
  U322
  (
    .A(n110),
    .B(n111),
    .Y(n447)
  );


  sky130_fd_sc_hd__xnor2_1
  U323
  (
    .A(A[15]),
    .B(n448),
    .Y(n110)
  );


  sky130_fd_sc_hd__o22ai_1
  U324
  (
    .A1(n107),
    .A2(n106),
    .B1(n449),
    .B2(n105),
    .Y(n111)
  );


  sky130_fd_sc_hd__and2_0
  U325
  (
    .A(n106),
    .B(n107),
    .X(n449)
  );


  sky130_fd_sc_hd__xnor2_1
  U326
  (
    .A(n97),
    .B(n450),
    .Y(n106)
  );


  sky130_fd_sc_hd__clkinv_1
  U327
  (
    .A(n413),
    .Y(n331)
  );


  sky130_fd_sc_hd__o22ai_1
  U328
  (
    .A1(n451),
    .A2(n452),
    .B1(n453),
    .B2(n454),
    .Y(n413)
  );


  sky130_fd_sc_hd__and2_0
  U329
  (
    .A(n452),
    .B(n451),
    .X(n453)
  );


  sky130_fd_sc_hd__clkinv_1
  U330
  (
    .A(n405),
    .Y(n351)
  );


  sky130_fd_sc_hd__o22ai_1
  U331
  (
    .A1(n455),
    .A2(n456),
    .B1(n457),
    .B2(n458),
    .Y(n405)
  );


  sky130_fd_sc_hd__and2_0
  U332
  (
    .A(n456),
    .B(n455),
    .X(n457)
  );


  sky130_fd_sc_hd__mux2i_1
  U333
  (
    .A0(n459),
    .A1(n460),
    .S(MODE_0_0),
    .Y(Y[0])
  );


  sky130_fd_sc_hd__xor2_1
  U334
  (
    .A(n461),
    .B(n462),
    .X(n460)
  );


  sky130_fd_sc_hd__xor2_1
  U335
  (
    .A(n463),
    .B(n464),
    .X(n462)
  );


  sky130_fd_sc_hd__maj3_1
  U336
  (
    .A(n465),
    .B(n164),
    .C(n466),
    .X(n464)
  );


  sky130_fd_sc_hd__maj3_1
  U337
  (
    .A(n467),
    .B(n171),
    .C(n468),
    .X(n466)
  );


  sky130_fd_sc_hd__a22oi_1
  U338
  (
    .A1(n469),
    .A2(n470),
    .B1(A[1]),
    .B2(n471),
    .Y(n468)
  );


  sky130_fd_sc_hd__maj3_1
  U339
  (
    .A(n472),
    .B(n473),
    .C(n474),
    .X(n467)
  );


  sky130_fd_sc_hd__a21oi_1
  U340
  (
    .A1(n475),
    .A2(n476),
    .B1(n477),
    .Y(n474)
  );


  sky130_fd_sc_hd__a22oi_1
  U341
  (
    .A1(n469),
    .A2(n478),
    .B1(n470),
    .B2(n471),
    .Y(n472)
  );


  sky130_fd_sc_hd__xnor2_1
  U342
  (
    .A(n479),
    .B(n480),
    .Y(n164)
  );


  sky130_fd_sc_hd__xor2_1
  U343
  (
    .A(n481),
    .B(n482),
    .X(n480)
  );


  sky130_fd_sc_hd__o21ai_0
  U344
  (
    .A1(n469),
    .A2(n471),
    .B1(A[1]),
    .Y(n479)
  );


  sky130_fd_sc_hd__maj3_1
  U345
  (
    .A(n483),
    .B(n115),
    .C(n484),
    .X(n465)
  );


  sky130_fd_sc_hd__maj3_1
  U346
  (
    .A(n485),
    .B(n229),
    .C(n486),
    .X(n484)
  );


  sky130_fd_sc_hd__a22oi_1
  U347
  (
    .A1(n487),
    .A2(B[3]),
    .B1(B[2]),
    .B2(n488),
    .Y(n486)
  );


  sky130_fd_sc_hd__maj3_1
  U348
  (
    .A(n489),
    .B(n490),
    .C(n491),
    .X(n485)
  );


  sky130_fd_sc_hd__a22oi_1
  U349
  (
    .A1(n469),
    .A2(n492),
    .B1(n478),
    .B2(n471),
    .Y(n491)
  );


  sky130_fd_sc_hd__a22oi_1
  U350
  (
    .A1(n493),
    .A2(n494),
    .B1(A[3]),
    .B2(n495),
    .Y(n489)
  );


  sky130_fd_sc_hd__xor2_1
  U351
  (
    .A(n169),
    .B(n496),
    .X(n115)
  );


  sky130_fd_sc_hd__xor2_1
  U352
  (
    .A(n171),
    .B(n168),
    .X(n496)
  );


  sky130_fd_sc_hd__o22ai_1
  U353
  (
    .A1(n497),
    .A2(n498),
    .B1(n499),
    .B2(n500),
    .Y(n168)
  );


  sky130_fd_sc_hd__o22ai_1
  U354
  (
    .A1(n501),
    .A2(n502),
    .B1(n473),
    .B2(n503),
    .Y(n169)
  );


  sky130_fd_sc_hd__nor2_1
  U355
  (
    .A(n504),
    .B(n505),
    .Y(n503)
  );


  sky130_fd_sc_hd__maj3_1
  U356
  (
    .A(n506),
    .B(n86),
    .C(n507),
    .X(n483)
  );


  sky130_fd_sc_hd__maj3_1
  U357
  (
    .A(n508),
    .B(n225),
    .C(n509),
    .X(n507)
  );


  sky130_fd_sc_hd__maj3_1
  U358
  (
    .A(n510),
    .B(n511),
    .C(n512),
    .X(n509)
  );


  sky130_fd_sc_hd__a21oi_1
  U359
  (
    .A1(n513),
    .A2(n514),
    .B1(n515),
    .Y(n512)
  );


  sky130_fd_sc_hd__a22oi_1
  U360
  (
    .A1(n469),
    .A2(n516),
    .B1(n492),
    .B2(n471),
    .Y(n510)
  );


  sky130_fd_sc_hd__maj3_1
  U361
  (
    .A(n517),
    .B(n518),
    .C(n519),
    .X(n508)
  );


  sky130_fd_sc_hd__a22oi_1
  U362
  (
    .A1(n493),
    .A2(n520),
    .B1(n494),
    .B2(n495),
    .Y(n519)
  );


  sky130_fd_sc_hd__maj3_1
  U363
  (
    .A(n521),
    .B(n522),
    .C(n523),
    .X(n517)
  );


  sky130_fd_sc_hd__a22oi_1
  U364
  (
    .A1(n487),
    .A2(B[6]),
    .B1(B[5]),
    .B2(n488),
    .Y(n523)
  );


  sky130_fd_sc_hd__a22oi_1
  U365
  (
    .A1(n469),
    .A2(n524),
    .B1(n516),
    .B2(n471),
    .Y(n521)
  );


  sky130_fd_sc_hd__xnor2_1
  U366
  (
    .A(n525),
    .B(n229),
    .Y(n86)
  );


  sky130_fd_sc_hd__xor2_1
  U367
  (
    .A(n502),
    .B(n526),
    .X(n229)
  );


  sky130_fd_sc_hd__xor2_1
  U368
  (
    .A(n473),
    .B(n501),
    .X(n526)
  );


  sky130_fd_sc_hd__clkinv_1
  U369
  (
    .A(n504),
    .Y(n501)
  );


  sky130_fd_sc_hd__o22ai_1
  U370
  (
    .A1(n497),
    .A2(n499),
    .B1(n527),
    .B2(n500),
    .Y(n504)
  );


  sky130_fd_sc_hd__clkinv_1
  U371
  (
    .A(n470),
    .Y(n499)
  );


  sky130_fd_sc_hd__xnor2_1
  U372
  (
    .A(n528),
    .B(A[1]),
    .Y(n470)
  );


  sky130_fd_sc_hd__clkinv_1
  U373
  (
    .A(n490),
    .Y(n473)
  );


  sky130_fd_sc_hd__clkinv_1
  U374
  (
    .A(n505),
    .Y(n502)
  );


  sky130_fd_sc_hd__o21ai_0
  U375
  (
    .A1(n493),
    .A2(n495),
    .B1(A[3]),
    .Y(n505)
  );


  sky130_fd_sc_hd__xnor2_1
  U376
  (
    .A(n227),
    .B(n226),
    .Y(n525)
  );


  sky130_fd_sc_hd__o22ai_1
  U377
  (
    .A1(n529),
    .A2(n530),
    .B1(n531),
    .B2(n532),
    .Y(n226)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U378
  (
    .B1(n533),
    .B2(n490),
    .A1_N(n534),
    .A2_N(n535),
    .Y(n227)
  );


  sky130_fd_sc_hd__nor2_1
  U379
  (
    .A(n534),
    .B(n535),
    .Y(n533)
  );


  sky130_fd_sc_hd__maj3_1
  U380
  (
    .A(n536),
    .B(n77),
    .C(n537),
    .X(n506)
  );


  sky130_fd_sc_hd__maj3_1
  U381
  (
    .A(n538),
    .B(n221),
    .C(n539),
    .X(n537)
  );


  sky130_fd_sc_hd__xor2_1
  U382
  (
    .A(n540),
    .B(n541),
    .X(n539)
  );


  sky130_fd_sc_hd__xor2_1
  U383
  (
    .A(n542),
    .B(n543),
    .X(n541)
  );


  sky130_fd_sc_hd__maj3_1
  U384
  (
    .A(n544),
    .B(n545),
    .C(n546),
    .X(n538)
  );


  sky130_fd_sc_hd__a22oi_1
  U385
  (
    .A1(n493),
    .A2(n547),
    .B1(n520),
    .B2(n495),
    .Y(n546)
  );


  sky130_fd_sc_hd__maj3_1
  U386
  (
    .A(n548),
    .B(n522),
    .C(n549),
    .X(n544)
  );


  sky130_fd_sc_hd__a22oi_1
  U387
  (
    .A1(n469),
    .A2(n550),
    .B1(n524),
    .B2(n471),
    .Y(n549)
  );


  sky130_fd_sc_hd__a22oi_1
  U388
  (
    .A1(n493),
    .A2(n551),
    .B1(n547),
    .B2(n495),
    .Y(n548)
  );


  sky130_fd_sc_hd__xnor2_1
  U389
  (
    .A(n552),
    .B(n225),
    .Y(n77)
  );


  sky130_fd_sc_hd__xor2_1
  U390
  (
    .A(n535),
    .B(n553),
    .X(n225)
  );


  sky130_fd_sc_hd__xor2_1
  U391
  (
    .A(n490),
    .B(n534),
    .X(n553)
  );


  sky130_fd_sc_hd__o22ai_1
  U392
  (
    .A1(n475),
    .A2(n477),
    .B1(n554),
    .B2(n476),
    .Y(n534)
  );


  sky130_fd_sc_hd__o22ai_1
  U393
  (
    .A1(n529),
    .A2(n531),
    .B1(n555),
    .B2(n532),
    .Y(n490)
  );


  sky130_fd_sc_hd__o22ai_1
  U394
  (
    .A1(n497),
    .A2(n527),
    .B1(n556),
    .B2(n500),
    .Y(n535)
  );


  sky130_fd_sc_hd__clkinv_1
  U395
  (
    .A(n478),
    .Y(n527)
  );


  sky130_fd_sc_hd__xnor2_1
  U396
  (
    .A(n557),
    .B(A[1]),
    .Y(n478)
  );


  sky130_fd_sc_hd__xnor2_1
  U397
  (
    .A(n223),
    .B(n222),
    .Y(n552)
  );


  sky130_fd_sc_hd__o22ai_1
  U398
  (
    .A1(n558),
    .A2(n559),
    .B1(n511),
    .B2(n560),
    .Y(n222)
  );


  sky130_fd_sc_hd__nor2_1
  U399
  (
    .A(n561),
    .B(n562),
    .Y(n560)
  );


  sky130_fd_sc_hd__o22ai_1
  U400
  (
    .A1(n543),
    .A2(n563),
    .B1(n518),
    .B2(n564),
    .Y(n223)
  );


  sky130_fd_sc_hd__nor2_1
  U401
  (
    .A(n565),
    .B(n540),
    .Y(n564)
  );


  sky130_fd_sc_hd__clkinv_1
  U402
  (
    .A(n540),
    .Y(n563)
  );


  sky130_fd_sc_hd__maj3_1
  U403
  (
    .A(n566),
    .B(n66),
    .C(n567),
    .X(n536)
  );


  sky130_fd_sc_hd__maj3_1
  U404
  (
    .A(n568),
    .B(n217),
    .C(n569),
    .X(n567)
  );


  sky130_fd_sc_hd__xor2_1
  U405
  (
    .A(n570),
    .B(n571),
    .X(n569)
  );


  sky130_fd_sc_hd__xor2_1
  U406
  (
    .A(n572),
    .B(n545),
    .X(n571)
  );


  sky130_fd_sc_hd__maj3_1
  U407
  (
    .A(n573),
    .B(A[7]),
    .C(n574),
    .X(n568)
  );


  sky130_fd_sc_hd__maj3_1
  U408
  (
    .A(n575),
    .B(n576),
    .C(n577),
    .X(n573)
  );


  sky130_fd_sc_hd__a22oi_1
  U409
  (
    .A1(n469),
    .A2(n578),
    .B1(n550),
    .B2(n471),
    .Y(n577)
  );


  sky130_fd_sc_hd__a22oi_1
  U410
  (
    .A1(n579),
    .A2(n580),
    .B1(n581),
    .B2(n582),
    .Y(n575)
  );


  sky130_fd_sc_hd__xnor2_1
  U411
  (
    .A(n583),
    .B(n221),
    .Y(n66)
  );


  sky130_fd_sc_hd__xor2_1
  U412
  (
    .A(n559),
    .B(n584),
    .X(n221)
  );


  sky130_fd_sc_hd__xor2_1
  U413
  (
    .A(n511),
    .B(n558),
    .X(n584)
  );


  sky130_fd_sc_hd__clkinv_1
  U414
  (
    .A(n561),
    .Y(n558)
  );


  sky130_fd_sc_hd__o22ai_1
  U415
  (
    .A1(n497),
    .A2(n556),
    .B1(n585),
    .B2(n500),
    .Y(n561)
  );


  sky130_fd_sc_hd__clkinv_1
  U416
  (
    .A(n492),
    .Y(n556)
  );


  sky130_fd_sc_hd__xnor2_1
  U417
  (
    .A(n530),
    .B(A[1]),
    .Y(n492)
  );


  sky130_fd_sc_hd__clkinv_1
  U418
  (
    .A(n562),
    .Y(n559)
  );


  sky130_fd_sc_hd__o21ai_0
  U419
  (
    .A1(n579),
    .A2(n582),
    .B1(A[5]),
    .Y(n562)
  );


  sky130_fd_sc_hd__xnor2_1
  U420
  (
    .A(n218),
    .B(n219),
    .Y(n583)
  );


  sky130_fd_sc_hd__xnor2_1
  U421
  (
    .A(n540),
    .B(n586),
    .Y(n219)
  );


  sky130_fd_sc_hd__xor2_1
  U422
  (
    .A(n518),
    .B(n543),
    .X(n586)
  );


  sky130_fd_sc_hd__clkinv_1
  U423
  (
    .A(n565),
    .Y(n543)
  );


  sky130_fd_sc_hd__o22ai_1
  U424
  (
    .A1(n475),
    .A2(n554),
    .B1(n587),
    .B2(n476),
    .Y(n565)
  );


  sky130_fd_sc_hd__clkinv_1
  U425
  (
    .A(n494),
    .Y(n554)
  );


  sky130_fd_sc_hd__xnor2_1
  U426
  (
    .A(n528),
    .B(A[3]),
    .Y(n494)
  );


  sky130_fd_sc_hd__clkinv_1
  U427
  (
    .A(n542),
    .Y(n518)
  );


  sky130_fd_sc_hd__o22ai_1
  U428
  (
    .A1(n529),
    .A2(n555),
    .B1(n588),
    .B2(n532),
    .Y(n542)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U429
  (
    .B1(n589),
    .B2(n522),
    .A1_N(n590),
    .A2_N(n591),
    .Y(n540)
  );


  sky130_fd_sc_hd__nor2_1
  U430
  (
    .A(n590),
    .B(n591),
    .Y(n589)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U431
  (
    .B1(n572),
    .B2(n570),
    .A1_N(n545),
    .A2_N(n592),
    .Y(n218)
  );


  sky130_fd_sc_hd__nor2_1
  U432
  (
    .A(n572),
    .B(n570),
    .Y(n592)
  );


  sky130_fd_sc_hd__maj3_1
  U433
  (
    .A(n593),
    .B(n57),
    .C(n594),
    .X(n566)
  );


  sky130_fd_sc_hd__maj3_1
  U434
  (
    .A(n595),
    .B(n213),
    .C(n596),
    .X(n594)
  );


  sky130_fd_sc_hd__xor2_1
  U435
  (
    .A(n597),
    .B(n598),
    .X(n596)
  );


  sky130_fd_sc_hd__xor2_1
  U436
  (
    .A(n599),
    .B(n574),
    .X(n598)
  );


  sky130_fd_sc_hd__maj3_1
  U437
  (
    .A(n600),
    .B(n601),
    .C(n602),
    .X(n595)
  );


  sky130_fd_sc_hd__a22oi_1
  U438
  (
    .A1(n493),
    .A2(n603),
    .B1(n551),
    .B2(n495),
    .Y(n602)
  );


  sky130_fd_sc_hd__maj3_1
  U439
  (
    .A(n604),
    .B(n605),
    .C(n606),
    .X(n600)
  );


  sky130_fd_sc_hd__a22oi_1
  U440
  (
    .A1(n607),
    .A2(n608),
    .B1(A[8]),
    .B2(n609),
    .Y(n606)
  );


  sky130_fd_sc_hd__a22oi_1
  U441
  (
    .A1(n469),
    .A2(n610),
    .B1(n578),
    .B2(n471),
    .Y(n604)
  );


  sky130_fd_sc_hd__xnor2_1
  U442
  (
    .A(n611),
    .B(n217),
    .Y(n57)
  );


  sky130_fd_sc_hd__xnor2_1
  U443
  (
    .A(n612),
    .B(n591),
    .Y(n217)
  );


  sky130_fd_sc_hd__o22ai_1
  U444
  (
    .A1(n497),
    .A2(n585),
    .B1(n613),
    .B2(n500),
    .Y(n591)
  );


  sky130_fd_sc_hd__clkinv_1
  U445
  (
    .A(n516),
    .Y(n585)
  );


  sky130_fd_sc_hd__xnor2_1
  U446
  (
    .A(n531),
    .B(A[1]),
    .Y(n516)
  );


  sky130_fd_sc_hd__xor2_1
  U447
  (
    .A(n590),
    .B(n511),
    .X(n612)
  );


  sky130_fd_sc_hd__clkinv_1
  U448
  (
    .A(n522),
    .Y(n511)
  );


  sky130_fd_sc_hd__o22ai_1
  U449
  (
    .A1(n529),
    .A2(n588),
    .B1(n614),
    .B2(n532),
    .Y(n590)
  );


  sky130_fd_sc_hd__xnor2_1
  U450
  (
    .A(n214),
    .B(n215),
    .Y(n611)
  );


  sky130_fd_sc_hd__xnor2_1
  U451
  (
    .A(n570),
    .B(n615),
    .Y(n215)
  );


  sky130_fd_sc_hd__xnor2_1
  U452
  (
    .A(n545),
    .B(n572),
    .Y(n615)
  );


  sky130_fd_sc_hd__o22ai_1
  U453
  (
    .A1(n475),
    .A2(n587),
    .B1(n616),
    .B2(n476),
    .Y(n572)
  );


  sky130_fd_sc_hd__clkinv_1
  U454
  (
    .A(n520),
    .Y(n587)
  );


  sky130_fd_sc_hd__xnor2_1
  U455
  (
    .A(n557),
    .B(A[3]),
    .Y(n520)
  );


  sky130_fd_sc_hd__a22oi_1
  U456
  (
    .A1(n582),
    .A2(A[5]),
    .B1(n617),
    .B2(n579),
    .Y(n545)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U457
  (
    .B1(n618),
    .B2(n522),
    .A1_N(n619),
    .A2_N(n620),
    .Y(n570)
  );


  sky130_fd_sc_hd__nor2_1
  U458
  (
    .A(n619),
    .B(n620),
    .Y(n618)
  );


  sky130_fd_sc_hd__o22a_1
  U459
  (
    .A1(n574),
    .A2(n621),
    .B1(A[7]),
    .B2(n622),
    .X(n214)
  );


  sky130_fd_sc_hd__and2_0
  U460
  (
    .A(n574),
    .B(n621),
    .X(n622)
  );


  sky130_fd_sc_hd__clkinv_1
  U461
  (
    .A(n597),
    .Y(n621)
  );


  sky130_fd_sc_hd__maj3_1
  U462
  (
    .A(n623),
    .B(n47),
    .C(n624),
    .X(n593)
  );


  sky130_fd_sc_hd__maj3_1
  U463
  (
    .A(n625),
    .B(n209),
    .C(n626),
    .X(n624)
  );


  sky130_fd_sc_hd__a21oi_1
  U464
  (
    .A1(n627),
    .A2(n628),
    .B1(n629),
    .Y(n626)
  );


  sky130_fd_sc_hd__a21oi_1
  U465
  (
    .A1(n630),
    .A2(n631),
    .B1(n632),
    .Y(n629)
  );


  sky130_fd_sc_hd__xor2_1
  U466
  (
    .A(n633),
    .B(n634),
    .X(n625)
  );


  sky130_fd_sc_hd__xor2_1
  U467
  (
    .A(n635),
    .B(n636),
    .X(n634)
  );


  sky130_fd_sc_hd__xnor2_1
  U468
  (
    .A(n637),
    .B(n213),
    .Y(n47)
  );


  sky130_fd_sc_hd__xor2_1
  U469
  (
    .A(n620),
    .B(n638),
    .X(n213)
  );


  sky130_fd_sc_hd__xor2_1
  U470
  (
    .A(n522),
    .B(n619),
    .X(n638)
  );


  sky130_fd_sc_hd__o22ai_1
  U471
  (
    .A1(n475),
    .A2(n616),
    .B1(n639),
    .B2(n476),
    .Y(n619)
  );


  sky130_fd_sc_hd__clkinv_1
  U472
  (
    .A(n547),
    .Y(n616)
  );


  sky130_fd_sc_hd__xnor2_1
  U473
  (
    .A(n530),
    .B(A[3]),
    .Y(n547)
  );


  sky130_fd_sc_hd__o22ai_1
  U474
  (
    .A1(n529),
    .A2(n614),
    .B1(n640),
    .B2(n532),
    .Y(n522)
  );


  sky130_fd_sc_hd__o22ai_1
  U475
  (
    .A1(n497),
    .A2(n613),
    .B1(n641),
    .B2(n500),
    .Y(n620)
  );


  sky130_fd_sc_hd__clkinv_1
  U476
  (
    .A(n524),
    .Y(n613)
  );


  sky130_fd_sc_hd__xnor2_1
  U477
  (
    .A(n555),
    .B(A[1]),
    .Y(n524)
  );


  sky130_fd_sc_hd__xnor2_1
  U478
  (
    .A(n210),
    .B(n211),
    .Y(n637)
  );


  sky130_fd_sc_hd__xnor2_1
  U479
  (
    .A(n597),
    .B(n642),
    .Y(n211)
  );


  sky130_fd_sc_hd__xor2_1
  U480
  (
    .A(A[7]),
    .B(n574),
    .X(n642)
  );


  sky130_fd_sc_hd__a22oi_1
  U481
  (
    .A1(n579),
    .A2(n581),
    .B1(n617),
    .B2(n582),
    .Y(n574)
  );


  sky130_fd_sc_hd__xnor2_1
  U482
  (
    .A(n528),
    .B(A[5]),
    .Y(n617)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U483
  (
    .B1(n576),
    .B2(n643),
    .A1_N(n644),
    .A2_N(n645),
    .Y(n597)
  );


  sky130_fd_sc_hd__nor2_1
  U484
  (
    .A(n644),
    .B(n645),
    .Y(n643)
  );


  sky130_fd_sc_hd__o22a_1
  U485
  (
    .A1(n636),
    .A2(n646),
    .B1(n601),
    .B2(n647),
    .X(n210)
  );


  sky130_fd_sc_hd__nor2_1
  U486
  (
    .A(n648),
    .B(n633),
    .Y(n647)
  );


  sky130_fd_sc_hd__clkinv_1
  U487
  (
    .A(n633),
    .Y(n646)
  );


  sky130_fd_sc_hd__maj3_1
  U488
  (
    .A(n649),
    .B(n36),
    .C(n650),
    .X(n623)
  );


  sky130_fd_sc_hd__a21oi_1
  U489
  (
    .A1(n205),
    .A2(n204),
    .B1(n651),
    .Y(n650)
  );


  sky130_fd_sc_hd__a21oi_1
  U490
  (
    .A1(n201),
    .A2(n200),
    .B1(n203),
    .Y(n651)
  );


  sky130_fd_sc_hd__clkinv_1
  U491
  (
    .A(n201),
    .Y(n205)
  );


  sky130_fd_sc_hd__xnor2_1
  U492
  (
    .A(n652),
    .B(n209),
    .Y(n36)
  );


  sky130_fd_sc_hd__xnor2_1
  U493
  (
    .A(n645),
    .B(n653),
    .Y(n209)
  );


  sky130_fd_sc_hd__xnor2_1
  U494
  (
    .A(n576),
    .B(n644),
    .Y(n653)
  );


  sky130_fd_sc_hd__a22o_1
  U495
  (
    .A1(n582),
    .A2(n581),
    .B1(n580),
    .B2(n579),
    .X(n644)
  );


  sky130_fd_sc_hd__xor2_1
  U496
  (
    .A(n557),
    .B(n515),
    .X(n581)
  );


  sky130_fd_sc_hd__a22oi_1
  U497
  (
    .A1(n488),
    .A2(B[7]),
    .B1(B[8]),
    .B2(n487),
    .Y(n576)
  );


  sky130_fd_sc_hd__o22ai_1
  U498
  (
    .A1(n497),
    .A2(n641),
    .B1(n654),
    .B2(n500),
    .Y(n645)
  );


  sky130_fd_sc_hd__clkinv_1
  U499
  (
    .A(n550),
    .Y(n641)
  );


  sky130_fd_sc_hd__xnor2_1
  U500
  (
    .A(n588),
    .B(A[1]),
    .Y(n550)
  );


  sky130_fd_sc_hd__xnor2_1
  U501
  (
    .A(n207),
    .B(n206),
    .Y(n652)
  );


  sky130_fd_sc_hd__o22a_1
  U502
  (
    .A1(n630),
    .A2(n631),
    .B1(n632),
    .B2(n655),
    .X(n206)
  );


  sky130_fd_sc_hd__nor2_1
  U503
  (
    .A(n627),
    .B(n628),
    .Y(n655)
  );


  sky130_fd_sc_hd__clkinv_1
  U504
  (
    .A(n628),
    .Y(n630)
  );


  sky130_fd_sc_hd__xnor2_1
  U505
  (
    .A(n633),
    .B(n656),
    .Y(n207)
  );


  sky130_fd_sc_hd__xor2_1
  U506
  (
    .A(n601),
    .B(n636),
    .X(n656)
  );


  sky130_fd_sc_hd__clkinv_1
  U507
  (
    .A(n648),
    .Y(n636)
  );


  sky130_fd_sc_hd__o22ai_1
  U508
  (
    .A1(n475),
    .A2(n639),
    .B1(n657),
    .B2(n476),
    .Y(n648)
  );


  sky130_fd_sc_hd__clkinv_1
  U509
  (
    .A(n551),
    .Y(n639)
  );


  sky130_fd_sc_hd__xnor2_1
  U510
  (
    .A(n531),
    .B(A[3]),
    .Y(n551)
  );


  sky130_fd_sc_hd__clkinv_1
  U511
  (
    .A(n635),
    .Y(n601)
  );


  sky130_fd_sc_hd__o22ai_1
  U512
  (
    .A1(n599),
    .A2(n301),
    .B1(n658),
    .B2(n659),
    .Y(n635)
  );


  sky130_fd_sc_hd__clkinv_1
  U513
  (
    .A(A[7]),
    .Y(n599)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U514
  (
    .B1(n660),
    .B2(n605),
    .A1_N(n661),
    .A2_N(n662),
    .Y(n633)
  );


  sky130_fd_sc_hd__nor2_1
  U515
  (
    .A(n661),
    .B(n662),
    .Y(n660)
  );


  sky130_fd_sc_hd__maj3_1
  U516
  (
    .A(n663),
    .B(n26),
    .C(n664),
    .X(n649)
  );


  sky130_fd_sc_hd__a21oi_1
  U517
  (
    .A1(n198),
    .A2(n199),
    .B1(n665),
    .Y(n664)
  );


  sky130_fd_sc_hd__a21oi_1
  U518
  (
    .A1(n194),
    .A2(n195),
    .B1(n197),
    .Y(n665)
  );


  sky130_fd_sc_hd__clkinv_1
  U519
  (
    .A(n194),
    .Y(n199)
  );


  sky130_fd_sc_hd__clkinv_1
  U520
  (
    .A(n195),
    .Y(n198)
  );


  sky130_fd_sc_hd__xor2_1
  U521
  (
    .A(n666),
    .B(n203),
    .X(n26)
  );


  sky130_fd_sc_hd__xnor2_1
  U522
  (
    .A(n667),
    .B(n662),
    .Y(n203)
  );


  sky130_fd_sc_hd__o22ai_1
  U523
  (
    .A1(n497),
    .A2(n654),
    .B1(n668),
    .B2(n500),
    .Y(n662)
  );


  sky130_fd_sc_hd__clkinv_1
  U524
  (
    .A(n578),
    .Y(n654)
  );


  sky130_fd_sc_hd__xnor2_1
  U525
  (
    .A(n614),
    .B(A[1]),
    .Y(n578)
  );


  sky130_fd_sc_hd__xnor2_1
  U526
  (
    .A(n661),
    .B(n605),
    .Y(n667)
  );


  sky130_fd_sc_hd__nand2_1
  U527
  (
    .A(B[8]),
    .B(n488),
    .Y(n605)
  );


  sky130_fd_sc_hd__o22ai_1
  U528
  (
    .A1(n658),
    .A2(n301),
    .B1(n669),
    .B2(n659),
    .Y(n661)
  );


  sky130_fd_sc_hd__clkinv_1
  U529
  (
    .A(n609),
    .Y(n658)
  );


  sky130_fd_sc_hd__xnor2_1
  U530
  (
    .A(n528),
    .B(A[7]),
    .Y(n609)
  );


  sky130_fd_sc_hd__xor2_1
  U531
  (
    .A(n201),
    .B(n200),
    .X(n666)
  );


  sky130_fd_sc_hd__clkinv_1
  U532
  (
    .A(n204),
    .Y(n200)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U533
  (
    .B1(n670),
    .B2(n671),
    .A1_N(n672),
    .A2_N(n673),
    .Y(n204)
  );


  sky130_fd_sc_hd__nor2_1
  U534
  (
    .A(n673),
    .B(n672),
    .Y(n670)
  );


  sky130_fd_sc_hd__xor2_1
  U535
  (
    .A(n628),
    .B(n674),
    .X(n201)
  );


  sky130_fd_sc_hd__xor2_1
  U536
  (
    .A(n627),
    .B(n632),
    .X(n674)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U537
  (
    .B1(n582),
    .B2(n580),
    .A1_N(n675),
    .A2_N(n514),
    .Y(n632)
  );


  sky130_fd_sc_hd__xnor2_1
  U538
  (
    .A(n530),
    .B(A[5]),
    .Y(n580)
  );


  sky130_fd_sc_hd__clkinv_1
  U539
  (
    .A(n631),
    .Y(n627)
  );


  sky130_fd_sc_hd__nand2_1
  U540
  (
    .A(n676),
    .B(n677),
    .Y(n631)
  );


  sky130_fd_sc_hd__o22ai_1
  U541
  (
    .A1(n475),
    .A2(n657),
    .B1(n678),
    .B2(n476),
    .Y(n628)
  );


  sky130_fd_sc_hd__clkinv_1
  U542
  (
    .A(n603),
    .Y(n657)
  );


  sky130_fd_sc_hd__xnor2_1
  U543
  (
    .A(n555),
    .B(A[3]),
    .Y(n603)
  );


  sky130_fd_sc_hd__maj3_1
  U544
  (
    .A(n679),
    .B(n191),
    .C(n680),
    .X(n663)
  );


  sky130_fd_sc_hd__a21oi_1
  U545
  (
    .A1(n373),
    .A2(n374),
    .B1(n681),
    .Y(n680)
  );


  sky130_fd_sc_hd__a21oi_1
  U546
  (
    .A1(n369),
    .A2(n370),
    .B1(n372),
    .Y(n681)
  );


  sky130_fd_sc_hd__xor2_1
  U547
  (
    .A(n682),
    .B(n197),
    .X(n191)
  );


  sky130_fd_sc_hd__xnor2_1
  U548
  (
    .A(n677),
    .B(n676),
    .Y(n197)
  );


  sky130_fd_sc_hd__o22ai_1
  U549
  (
    .A1(n475),
    .A2(n678),
    .B1(n683),
    .B2(n476),
    .Y(n676)
  );


  sky130_fd_sc_hd__xor2_1
  U550
  (
    .A(n588),
    .B(A[3]),
    .X(n678)
  );


  sky130_fd_sc_hd__o22ai_1
  U551
  (
    .A1(n669),
    .A2(n301),
    .B1(n684),
    .B2(n659),
    .Y(n677)
  );


  sky130_fd_sc_hd__clkinv_1
  U552
  (
    .A(n608),
    .Y(n669)
  );


  sky130_fd_sc_hd__xnor2_1
  U553
  (
    .A(n557),
    .B(A[7]),
    .Y(n608)
  );


  sky130_fd_sc_hd__xor2_1
  U554
  (
    .A(n195),
    .B(n194),
    .X(n682)
  );


  sky130_fd_sc_hd__a22oi_1
  U555
  (
    .A1(n685),
    .A2(n686),
    .B1(n687),
    .B2(n688),
    .Y(n194)
  );


  sky130_fd_sc_hd__or2_0
  U556
  (
    .A(n686),
    .B(n685),
    .X(n687)
  );


  sky130_fd_sc_hd__xor2_1
  U557
  (
    .A(n673),
    .B(n689),
    .X(n195)
  );


  sky130_fd_sc_hd__xor2_1
  U558
  (
    .A(n671),
    .B(n672),
    .X(n689)
  );


  sky130_fd_sc_hd__o22ai_1
  U559
  (
    .A1(n497),
    .A2(n668),
    .B1(n690),
    .B2(n500),
    .Y(n672)
  );


  sky130_fd_sc_hd__xor2_1
  U560
  (
    .A(n498),
    .B(B[8]),
    .X(n690)
  );


  sky130_fd_sc_hd__clkinv_1
  U561
  (
    .A(n610),
    .Y(n668)
  );


  sky130_fd_sc_hd__xnor2_1
  U562
  (
    .A(n640),
    .B(A[1]),
    .Y(n610)
  );


  sky130_fd_sc_hd__o21ai_0
  U563
  (
    .A1(n691),
    .A2(n469),
    .B1(A[1]),
    .Y(n671)
  );


  sky130_fd_sc_hd__clkinv_1
  U564
  (
    .A(n500),
    .Y(n469)
  );


  sky130_fd_sc_hd__nor2_1
  U565
  (
    .A(B[8]),
    .B(n497),
    .Y(n691)
  );


  sky130_fd_sc_hd__o22ai_1
  U566
  (
    .A1(n513),
    .A2(n675),
    .B1(n692),
    .B2(n514),
    .Y(n673)
  );


  sky130_fd_sc_hd__xor2_1
  U567
  (
    .A(n531),
    .B(A[5]),
    .X(n675)
  );


  sky130_fd_sc_hd__maj3_1
  U568
  (
    .A(n693),
    .B(n358),
    .C(n694),
    .X(n679)
  );


  sky130_fd_sc_hd__a21oi_1
  U569
  (
    .A1(n380),
    .A2(n381),
    .B1(n695),
    .Y(n694)
  );


  sky130_fd_sc_hd__a21oi_1
  U570
  (
    .A1(n376),
    .A2(n377),
    .B1(n379),
    .Y(n695)
  );


  sky130_fd_sc_hd__xnor2_1
  U571
  (
    .A(n372),
    .B(n696),
    .Y(n358)
  );


  sky130_fd_sc_hd__xor2_1
  U572
  (
    .A(n373),
    .B(n369),
    .X(n696)
  );


  sky130_fd_sc_hd__clkinv_1
  U573
  (
    .A(n374),
    .Y(n369)
  );


  sky130_fd_sc_hd__o22ai_1
  U574
  (
    .A1(n513),
    .A2(n692),
    .B1(n697),
    .B2(n514),
    .Y(n374)
  );


  sky130_fd_sc_hd__xor2_1
  U575
  (
    .A(n555),
    .B(A[5]),
    .X(n692)
  );


  sky130_fd_sc_hd__clkinv_1
  U576
  (
    .A(n370),
    .Y(n373)
  );


  sky130_fd_sc_hd__nand2_1
  U577
  (
    .A(n698),
    .B(n699),
    .Y(n370)
  );


  sky130_fd_sc_hd__xnor2_1
  U578
  (
    .A(n700),
    .B(n686),
    .Y(n372)
  );


  sky130_fd_sc_hd__o22ai_1
  U579
  (
    .A1(n475),
    .A2(n683),
    .B1(n701),
    .B2(n476),
    .Y(n686)
  );


  sky130_fd_sc_hd__xor2_1
  U580
  (
    .A(n614),
    .B(A[3]),
    .X(n683)
  );


  sky130_fd_sc_hd__xor2_1
  U581
  (
    .A(n685),
    .B(n688),
    .X(n700)
  );


  sky130_fd_sc_hd__nor2_1
  U582
  (
    .A(n302),
    .B(n497),
    .Y(n688)
  );


  sky130_fd_sc_hd__o22ai_1
  U583
  (
    .A1(n684),
    .A2(n301),
    .B1(n702),
    .B2(n659),
    .Y(n685)
  );


  sky130_fd_sc_hd__xor2_1
  U584
  (
    .A(n530),
    .B(A[7]),
    .X(n684)
  );


  sky130_fd_sc_hd__maj3_1
  U585
  (
    .A(n703),
    .B(n352),
    .C(n704),
    .X(n693)
  );


  sky130_fd_sc_hd__maj3_1
  U586
  (
    .A(n705),
    .B(n390),
    .C(n706),
    .X(n704)
  );


  sky130_fd_sc_hd__a22oi_1
  U587
  (
    .A1(n607),
    .A2(n707),
    .B1(A[8]),
    .B2(n708),
    .Y(n706)
  );


  sky130_fd_sc_hd__a22oi_1
  U588
  (
    .A1(n579),
    .A2(n709),
    .B1(n710),
    .B2(n582),
    .Y(n705)
  );


  sky130_fd_sc_hd__xnor2_1
  U589
  (
    .A(n379),
    .B(n711),
    .Y(n352)
  );


  sky130_fd_sc_hd__xor2_1
  U590
  (
    .A(n380),
    .B(n376),
    .X(n711)
  );


  sky130_fd_sc_hd__clkinv_1
  U591
  (
    .A(n381),
    .Y(n376)
  );


  sky130_fd_sc_hd__o22ai_1
  U592
  (
    .A1(n513),
    .A2(n697),
    .B1(n712),
    .B2(n514),
    .Y(n381)
  );


  sky130_fd_sc_hd__xor2_1
  U593
  (
    .A(n588),
    .B(A[5]),
    .X(n697)
  );


  sky130_fd_sc_hd__clkinv_1
  U594
  (
    .A(n377),
    .Y(n380)
  );


  sky130_fd_sc_hd__o21ai_0
  U595
  (
    .A1(n713),
    .A2(n493),
    .B1(A[3]),
    .Y(n377)
  );


  sky130_fd_sc_hd__clkinv_1
  U596
  (
    .A(n476),
    .Y(n493)
  );


  sky130_fd_sc_hd__nor2_1
  U597
  (
    .A(B[8]),
    .B(n475),
    .Y(n713)
  );


  sky130_fd_sc_hd__xnor2_1
  U598
  (
    .A(n699),
    .B(n698),
    .Y(n379)
  );


  sky130_fd_sc_hd__o22ai_1
  U599
  (
    .A1(n475),
    .A2(n701),
    .B1(n714),
    .B2(n476),
    .Y(n698)
  );


  sky130_fd_sc_hd__nand2_1
  U600
  (
    .A(n475),
    .B(n715),
    .Y(n476)
  );


  sky130_fd_sc_hd__xor2_1
  U601
  (
    .A(A[4]),
    .B(A[3]),
    .X(n715)
  );


  sky130_fd_sc_hd__xor2_1
  U602
  (
    .A(n477),
    .B(B[8]),
    .X(n714)
  );


  sky130_fd_sc_hd__clkinv_1
  U603
  (
    .A(A[3]),
    .Y(n477)
  );


  sky130_fd_sc_hd__xor2_1
  U604
  (
    .A(n640),
    .B(A[3]),
    .X(n701)
  );


  sky130_fd_sc_hd__clkinv_1
  U605
  (
    .A(n495),
    .Y(n475)
  );


  sky130_fd_sc_hd__o22ai_1
  U606
  (
    .A1(n702),
    .A2(n301),
    .B1(n716),
    .B2(n659),
    .Y(n699)
  );


  sky130_fd_sc_hd__xor2_1
  U607
  (
    .A(n531),
    .B(A[7]),
    .X(n702)
  );


  sky130_fd_sc_hd__clkinv_1
  U608
  (
    .A(B[3]),
    .Y(n531)
  );


  sky130_fd_sc_hd__a21oi_1
  U609
  (
    .A1(n345),
    .A2(n344),
    .B1(n717),
    .Y(n703)
  );


  sky130_fd_sc_hd__a21oi_1
  U610
  (
    .A1(n384),
    .A2(n385),
    .B1(n342),
    .Y(n717)
  );


  sky130_fd_sc_hd__xnor2_1
  U611
  (
    .A(n718),
    .B(n388),
    .Y(n342)
  );


  sky130_fd_sc_hd__o22ai_1
  U612
  (
    .A1(n513),
    .A2(n712),
    .B1(n719),
    .B2(n514),
    .Y(n388)
  );


  sky130_fd_sc_hd__clkinv_1
  U613
  (
    .A(n710),
    .Y(n712)
  );


  sky130_fd_sc_hd__xnor2_1
  U614
  (
    .A(n614),
    .B(A[5]),
    .Y(n710)
  );


  sky130_fd_sc_hd__xnor2_1
  U615
  (
    .A(n387),
    .B(n390),
    .Y(n718)
  );


  sky130_fd_sc_hd__nand2_1
  U616
  (
    .A(B[8]),
    .B(n495),
    .Y(n390)
  );


  sky130_fd_sc_hd__xnor2_1
  U617
  (
    .A(n720),
    .B(A[5]),
    .Y(n495)
  );


  sky130_fd_sc_hd__o22ai_1
  U618
  (
    .A1(n716),
    .A2(n301),
    .B1(n721),
    .B2(n659),
    .Y(n387)
  );


  sky130_fd_sc_hd__clkinv_1
  U619
  (
    .A(n708),
    .Y(n716)
  );


  sky130_fd_sc_hd__xnor2_1
  U620
  (
    .A(n555),
    .B(A[7]),
    .Y(n708)
  );


  sky130_fd_sc_hd__clkinv_1
  U621
  (
    .A(B[4]),
    .Y(n555)
  );


  sky130_fd_sc_hd__clkinv_1
  U622
  (
    .A(n384),
    .Y(n344)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U623
  (
    .B1(n334),
    .B2(n335),
    .A1_N(n722),
    .A2_N(n332),
    .Y(n384)
  );


  sky130_fd_sc_hd__xnor2_1
  U624
  (
    .A(n723),
    .B(n724),
    .Y(n332)
  );


  sky130_fd_sc_hd__nor2_1
  U625
  (
    .A(n335),
    .B(n334),
    .Y(n722)
  );


  sky130_fd_sc_hd__o22ai_1
  U626
  (
    .A1(n323),
    .A2(n324),
    .B1(n323),
    .B2(n325),
    .Y(n335)
  );


  sky130_fd_sc_hd__nand2_1
  U627
  (
    .A(B[8]),
    .B(n582),
    .Y(n325)
  );


  sky130_fd_sc_hd__nand2b_1
  U628
  (
    .A_N(n315),
    .B(n314),
    .Y(n324)
  );


  sky130_fd_sc_hd__o22ai_1
  U629
  (
    .A1(B[8]),
    .A2(n659),
    .B1(n725),
    .B2(n301),
    .Y(n314)
  );


  sky130_fd_sc_hd__a21oi_1
  U630
  (
    .A1(n302),
    .A2(A[7]),
    .B1(n607),
    .Y(n315)
  );


  sky130_fd_sc_hd__clkinv_1
  U631
  (
    .A(n659),
    .Y(n607)
  );


  sky130_fd_sc_hd__clkinv_1
  U632
  (
    .A(B[8]),
    .Y(n302)
  );


  sky130_fd_sc_hd__o22a_1
  U633
  (
    .A1(n726),
    .A2(n301),
    .B1(n725),
    .B2(n659),
    .X(n323)
  );


  sky130_fd_sc_hd__xor2_1
  U634
  (
    .A(n640),
    .B(A[7]),
    .X(n725)
  );


  sky130_fd_sc_hd__o22ai_1
  U635
  (
    .A1(n513),
    .A2(n719),
    .B1(n727),
    .B2(n514),
    .Y(n334)
  );


  sky130_fd_sc_hd__xor2_1
  U636
  (
    .A(n515),
    .B(B[8]),
    .X(n727)
  );


  sky130_fd_sc_hd__clkinv_1
  U637
  (
    .A(n709),
    .Y(n719)
  );


  sky130_fd_sc_hd__xnor2_1
  U638
  (
    .A(n640),
    .B(A[5]),
    .Y(n709)
  );


  sky130_fd_sc_hd__clkinv_1
  U639
  (
    .A(B[7]),
    .Y(n640)
  );


  sky130_fd_sc_hd__clkinv_1
  U640
  (
    .A(n385),
    .Y(n345)
  );


  sky130_fd_sc_hd__nand2_1
  U641
  (
    .A(n724),
    .B(n723),
    .Y(n385)
  );


  sky130_fd_sc_hd__o22ai_1
  U642
  (
    .A1(n721),
    .A2(n301),
    .B1(n726),
    .B2(n659),
    .Y(n723)
  );


  sky130_fd_sc_hd__nand2_1
  U643
  (
    .A(A[7]),
    .B(n301),
    .Y(n659)
  );


  sky130_fd_sc_hd__xor2_1
  U644
  (
    .A(n614),
    .B(A[7]),
    .X(n726)
  );


  sky130_fd_sc_hd__clkinv_1
  U645
  (
    .A(B[6]),
    .Y(n614)
  );


  sky130_fd_sc_hd__clkinv_1
  U646
  (
    .A(n707),
    .Y(n721)
  );


  sky130_fd_sc_hd__xnor2_1
  U647
  (
    .A(n588),
    .B(A[7]),
    .Y(n707)
  );


  sky130_fd_sc_hd__clkinv_1
  U648
  (
    .A(B[5]),
    .Y(n588)
  );


  sky130_fd_sc_hd__o21a_1
  U649
  (
    .A1(n728),
    .A2(n579),
    .B1(A[5]),
    .X(n724)
  );


  sky130_fd_sc_hd__clkinv_1
  U650
  (
    .A(n514),
    .Y(n579)
  );


  sky130_fd_sc_hd__nand2_1
  U651
  (
    .A(n513),
    .B(n729),
    .Y(n514)
  );


  sky130_fd_sc_hd__xor2_1
  U652
  (
    .A(A[6]),
    .B(A[5]),
    .X(n729)
  );


  sky130_fd_sc_hd__nor2_1
  U653
  (
    .A(B[8]),
    .B(n513),
    .Y(n728)
  );


  sky130_fd_sc_hd__clkinv_1
  U654
  (
    .A(n582),
    .Y(n513)
  );


  sky130_fd_sc_hd__xnor2_1
  U655
  (
    .A(n730),
    .B(A[7]),
    .Y(n582)
  );


  sky130_fd_sc_hd__clkinv_1
  U656
  (
    .A(A[6]),
    .Y(n730)
  );


  sky130_fd_sc_hd__maj3_1
  U657
  (
    .A(n731),
    .B(n481),
    .C(n482),
    .X(n463)
  );


  sky130_fd_sc_hd__a22oi_1
  U658
  (
    .A1(n487),
    .A2(B[1]),
    .B1(B[0]),
    .B2(n488),
    .Y(n482)
  );


  sky130_fd_sc_hd__clkinv_1
  U659
  (
    .A(n532),
    .Y(n487)
  );


  sky130_fd_sc_hd__clkinv_1
  U660
  (
    .A(n171),
    .Y(n481)
  );


  sky130_fd_sc_hd__o22ai_1
  U661
  (
    .A1(n529),
    .A2(n557),
    .B1(n530),
    .B2(n532),
    .Y(n171)
  );


  sky130_fd_sc_hd__clkinv_1
  U662
  (
    .A(B[2]),
    .Y(n530)
  );


  sky130_fd_sc_hd__clkinv_1
  U663
  (
    .A(B[1]),
    .Y(n557)
  );


  sky130_fd_sc_hd__a21oi_1
  U664
  (
    .A1(n497),
    .A2(n500),
    .B1(n498),
    .Y(n731)
  );


  sky130_fd_sc_hd__nand2_1
  U665
  (
    .A(n497),
    .B(n732),
    .Y(n500)
  );


  sky130_fd_sc_hd__xor2_1
  U666
  (
    .A(A[2]),
    .B(A[1]),
    .X(n732)
  );


  sky130_fd_sc_hd__clkinv_1
  U667
  (
    .A(n471),
    .Y(n497)
  );


  sky130_fd_sc_hd__xnor2_1
  U668
  (
    .A(n733),
    .B(A[3]),
    .Y(n471)
  );


  sky130_fd_sc_hd__nor2_1
  U669
  (
    .A(n528),
    .B(n532),
    .Y(n461)
  );


  sky130_fd_sc_hd__nand2_1
  U670
  (
    .A(n529),
    .B(A[0]),
    .Y(n532)
  );


  sky130_fd_sc_hd__clkinv_1
  U671
  (
    .A(n488),
    .Y(n529)
  );


  sky130_fd_sc_hd__xnor2_1
  U672
  (
    .A(n734),
    .B(A[1]),
    .Y(n488)
  );


  sky130_fd_sc_hd__clkinv_1
  U673
  (
    .A(A[0]),
    .Y(n734)
  );


  sky130_fd_sc_hd__clkinv_1
  U674
  (
    .A(B[0]),
    .Y(n528)
  );


  sky130_fd_sc_hd__xor2_1
  U675
  (
    .A(n735),
    .B(n736),
    .X(n459)
  );


  sky130_fd_sc_hd__xor2_1
  U676
  (
    .A(n737),
    .B(n738),
    .X(n736)
  );


  sky130_fd_sc_hd__nor2_1
  U677
  (
    .A(n236),
    .B(n739),
    .Y(n738)
  );


  sky130_fd_sc_hd__nand2_1
  U678
  (
    .A(n740),
    .B(n741),
    .Y(n737)
  );


  sky130_fd_sc_hd__xnor2_1
  U679
  (
    .A(n742),
    .B(n743),
    .Y(n735)
  );


  sky130_fd_sc_hd__maj3_1
  U680
  (
    .A(n744),
    .B(n231),
    .C(n745),
    .X(n743)
  );


  sky130_fd_sc_hd__maj3_1
  U681
  (
    .A(n746),
    .B(n236),
    .C(n747),
    .X(n745)
  );


  sky130_fd_sc_hd__a21oi_1
  U682
  (
    .A1(n748),
    .A2(n749),
    .B1(n750),
    .Y(n747)
  );


  sky130_fd_sc_hd__o21a_1
  U683
  (
    .A1(n749),
    .A2(n748),
    .B1(n751),
    .X(n750)
  );


  sky130_fd_sc_hd__xor2_1
  U684
  (
    .A(n740),
    .B(n752),
    .X(n746)
  );


  sky130_fd_sc_hd__xor2_1
  U685
  (
    .A(n753),
    .B(n754),
    .X(n231)
  );


  sky130_fd_sc_hd__xor2_1
  U686
  (
    .A(n755),
    .B(n236),
    .X(n753)
  );


  sky130_fd_sc_hd__maj3_1
  U687
  (
    .A(n756),
    .B(n118),
    .C(n757),
    .X(n744)
  );


  sky130_fd_sc_hd__maj3_1
  U688
  (
    .A(n758),
    .B(n291),
    .C(n759),
    .X(n757)
  );


  sky130_fd_sc_hd__xor2_1
  U689
  (
    .A(n740),
    .B(n760),
    .X(n759)
  );


  sky130_fd_sc_hd__a21oi_1
  U690
  (
    .A1(n761),
    .A2(n762),
    .B1(n763),
    .Y(n758)
  );


  sky130_fd_sc_hd__a21oi_1
  U691
  (
    .A1(n764),
    .A2(n765),
    .B1(n749),
    .Y(n763)
  );


  sky130_fd_sc_hd__xor2_1
  U692
  (
    .A(n235),
    .B(n766),
    .X(n118)
  );


  sky130_fd_sc_hd__xor2_1
  U693
  (
    .A(n236),
    .B(n234),
    .X(n766)
  );


  sky130_fd_sc_hd__clkinv_1
  U694
  (
    .A(n238),
    .Y(n234)
  );


  sky130_fd_sc_hd__maj3_1
  U695
  (
    .A(n749),
    .B(n751),
    .C(n748),
    .X(n238)
  );


  sky130_fd_sc_hd__xnor2_1
  U696
  (
    .A(n739),
    .B(n752),
    .Y(n235)
  );


  sky130_fd_sc_hd__a222oi_1
  U697
  (
    .A1(n767),
    .A2(n768),
    .B1(n769),
    .B2(n741),
    .C1(n770),
    .C2(n771),
    .Y(n752)
  );


  sky130_fd_sc_hd__maj3_1
  U698
  (
    .A(n772),
    .B(n90),
    .C(n773),
    .X(n756)
  );


  sky130_fd_sc_hd__maj3_1
  U699
  (
    .A(n774),
    .B(n287),
    .C(n775),
    .X(n773)
  );


  sky130_fd_sc_hd__xor2_1
  U700
  (
    .A(n740),
    .B(n776),
    .X(n775)
  );


  sky130_fd_sc_hd__xor2_1
  U701
  (
    .A(n751),
    .B(n777),
    .X(n774)
  );


  sky130_fd_sc_hd__xnor2_1
  U702
  (
    .A(n778),
    .B(n291),
    .Y(n90)
  );


  sky130_fd_sc_hd__xor2_1
  U703
  (
    .A(n749),
    .B(n779),
    .X(n291)
  );


  sky130_fd_sc_hd__xor2_1
  U704
  (
    .A(n780),
    .B(n748),
    .X(n779)
  );


  sky130_fd_sc_hd__nor2_1
  U705
  (
    .A(n781),
    .B(n739),
    .Y(n748)
  );


  sky130_fd_sc_hd__xnor2_1
  U706
  (
    .A(n289),
    .B(n288),
    .Y(n778)
  );


  sky130_fd_sc_hd__o22a_1
  U707
  (
    .A1(n764),
    .A2(n765),
    .B1(n749),
    .B2(n782),
    .X(n288)
  );


  sky130_fd_sc_hd__nor2_1
  U708
  (
    .A(n761),
    .B(n762),
    .Y(n782)
  );


  sky130_fd_sc_hd__clkinv_1
  U709
  (
    .A(n762),
    .Y(n764)
  );


  sky130_fd_sc_hd__xnor2_1
  U710
  (
    .A(n739),
    .B(n760),
    .Y(n289)
  );


  sky130_fd_sc_hd__a221oi_1
  U711
  (
    .A1(n783),
    .A2(n741),
    .B1(n771),
    .B2(n784),
    .C1(n785),
    .Y(n760)
  );


  sky130_fd_sc_hd__o22ai_1
  U712
  (
    .A1(n786),
    .A2(n787),
    .B1(n788),
    .B2(n789),
    .Y(n785)
  );


  sky130_fd_sc_hd__maj3_1
  U713
  (
    .A(n790),
    .B(n81),
    .C(n791),
    .X(n772)
  );


  sky130_fd_sc_hd__maj3_1
  U714
  (
    .A(n792),
    .B(n283),
    .C(n793),
    .X(n791)
  );


  sky130_fd_sc_hd__maj3_1
  U715
  (
    .A(n794),
    .B(n795),
    .C(n796),
    .X(n793)
  );


  sky130_fd_sc_hd__a21oi_1
  U716
  (
    .A1(n797),
    .A2(n798),
    .B1(n799),
    .Y(n796)
  );


  sky130_fd_sc_hd__a21oi_1
  U717
  (
    .A1(n800),
    .A2(n801),
    .B1(n802),
    .Y(n799)
  );


  sky130_fd_sc_hd__xor2_1
  U718
  (
    .A(n740),
    .B(n803),
    .X(n794)
  );


  sky130_fd_sc_hd__xor2_1
  U719
  (
    .A(n780),
    .B(n804),
    .X(n792)
  );


  sky130_fd_sc_hd__xnor2_1
  U720
  (
    .A(n805),
    .B(n284),
    .Y(n81)
  );


  sky130_fd_sc_hd__xor2_1
  U721
  (
    .A(n739),
    .B(n776),
    .X(n284)
  );


  sky130_fd_sc_hd__a221oi_1
  U722
  (
    .A1(n806),
    .A2(n771),
    .B1(n767),
    .B2(n807),
    .C1(n808),
    .Y(n776)
  );


  sky130_fd_sc_hd__o22ai_1
  U723
  (
    .A1(n786),
    .A2(n789),
    .B1(n788),
    .B2(n809),
    .Y(n808)
  );


  sky130_fd_sc_hd__xnor2_1
  U724
  (
    .A(n287),
    .B(n285),
    .Y(n805)
  );


  sky130_fd_sc_hd__xnor2_1
  U725
  (
    .A(n777),
    .B(n751),
    .Y(n285)
  );


  sky130_fd_sc_hd__o22ai_1
  U726
  (
    .A1(n810),
    .A2(n811),
    .B1(n812),
    .B2(n813),
    .Y(n777)
  );


  sky130_fd_sc_hd__xor2_1
  U727
  (
    .A(n762),
    .B(n814),
    .X(n287)
  );


  sky130_fd_sc_hd__xor2_1
  U728
  (
    .A(n761),
    .B(n749),
    .X(n814)
  );


  sky130_fd_sc_hd__nor2_1
  U729
  (
    .A(n815),
    .B(n739),
    .Y(n749)
  );


  sky130_fd_sc_hd__o22ai_1
  U730
  (
    .A1(n816),
    .A2(n817),
    .B1(n761),
    .B2(n818),
    .Y(n762)
  );


  sky130_fd_sc_hd__nor2_1
  U731
  (
    .A(n819),
    .B(n820),
    .Y(n818)
  );


  sky130_fd_sc_hd__maj3_1
  U732
  (
    .A(n821),
    .B(n70),
    .C(n822),
    .X(n790)
  );


  sky130_fd_sc_hd__maj3_1
  U733
  (
    .A(n823),
    .B(n279),
    .C(n824),
    .X(n822)
  );


  sky130_fd_sc_hd__xor2_1
  U734
  (
    .A(n780),
    .B(n825),
    .X(n824)
  );


  sky130_fd_sc_hd__maj3_1
  U735
  (
    .A(n826),
    .B(n827),
    .C(n828),
    .X(n823)
  );


  sky130_fd_sc_hd__maj3_1
  U736
  (
    .A(n829),
    .B(n802),
    .C(n830),
    .X(n828)
  );


  sky130_fd_sc_hd__a21oi_1
  U737
  (
    .A1(n831),
    .A2(n832),
    .B1(n833),
    .Y(n830)
  );


  sky130_fd_sc_hd__o21a_1
  U738
  (
    .A1(n832),
    .A2(n831),
    .B1(n834),
    .X(n833)
  );


  sky130_fd_sc_hd__xor2_1
  U739
  (
    .A(n740),
    .B(n835),
    .X(n829)
  );


  sky130_fd_sc_hd__maj3_1
  U740
  (
    .A(n836),
    .B(n837),
    .C(n838),
    .X(n826)
  );


  sky130_fd_sc_hd__maj3_1
  U741
  (
    .A(n839),
    .B(n840),
    .C(n841),
    .X(n838)
  );


  sky130_fd_sc_hd__xor2_1
  U742
  (
    .A(n740),
    .B(n842),
    .X(n841)
  );


  sky130_fd_sc_hd__a21oi_1
  U743
  (
    .A1(n843),
    .A2(n844),
    .B1(n845),
    .Y(n839)
  );


  sky130_fd_sc_hd__a21oi_1
  U744
  (
    .A1(n846),
    .A2(n847),
    .B1(n832),
    .Y(n845)
  );


  sky130_fd_sc_hd__xor2_1
  U745
  (
    .A(n780),
    .B(n848),
    .X(n836)
  );


  sky130_fd_sc_hd__xnor2_1
  U746
  (
    .A(n849),
    .B(n283),
    .Y(n70)
  );


  sky130_fd_sc_hd__xor2_1
  U747
  (
    .A(n817),
    .B(n850),
    .X(n283)
  );


  sky130_fd_sc_hd__xor2_1
  U748
  (
    .A(n761),
    .B(n816),
    .X(n850)
  );


  sky130_fd_sc_hd__clkinv_1
  U749
  (
    .A(n820),
    .Y(n816)
  );


  sky130_fd_sc_hd__maj3_1
  U750
  (
    .A(n802),
    .B(n851),
    .C(n852),
    .X(n820)
  );


  sky130_fd_sc_hd__clkinv_1
  U751
  (
    .A(n765),
    .Y(n761)
  );


  sky130_fd_sc_hd__nand2_1
  U752
  (
    .A(n740),
    .B(n853),
    .Y(n765)
  );


  sky130_fd_sc_hd__clkinv_1
  U753
  (
    .A(n819),
    .Y(n817)
  );


  sky130_fd_sc_hd__xor2_1
  U754
  (
    .A(n739),
    .B(n854),
    .X(n819)
  );


  sky130_fd_sc_hd__a221oi_1
  U755
  (
    .A1(n769),
    .A2(n807),
    .B1(n855),
    .B2(n771),
    .C1(n856),
    .Y(n854)
  );


  sky130_fd_sc_hd__o22ai_1
  U756
  (
    .A1(n815),
    .A2(n787),
    .B1(n786),
    .B2(n809),
    .Y(n856)
  );


  sky130_fd_sc_hd__xnor2_1
  U757
  (
    .A(n281),
    .B(n280),
    .Y(n849)
  );


  sky130_fd_sc_hd__o22a_1
  U758
  (
    .A1(n857),
    .A2(n858),
    .B1(n859),
    .B2(n795),
    .X(n280)
  );


  sky130_fd_sc_hd__and2_0
  U759
  (
    .A(n858),
    .B(n857),
    .X(n859)
  );


  sky130_fd_sc_hd__xnor2_1
  U760
  (
    .A(n751),
    .B(n804),
    .Y(n281)
  );


  sky130_fd_sc_hd__a222oi_1
  U761
  (
    .A1(n860),
    .A2(n768),
    .B1(n861),
    .B2(n741),
    .C1(n770),
    .C2(n862),
    .Y(n804)
  );


  sky130_fd_sc_hd__maj3_1
  U762
  (
    .A(n863),
    .B(n60),
    .C(n864),
    .X(n821)
  );


  sky130_fd_sc_hd__maj3_1
  U763
  (
    .A(n865),
    .B(n275),
    .C(n866),
    .X(n864)
  );


  sky130_fd_sc_hd__xor2_1
  U764
  (
    .A(n851),
    .B(n867),
    .X(n866)
  );


  sky130_fd_sc_hd__xor2_1
  U765
  (
    .A(n780),
    .B(n868),
    .X(n865)
  );


  sky130_fd_sc_hd__xnor2_1
  U766
  (
    .A(n869),
    .B(n279),
    .Y(n60)
  );


  sky130_fd_sc_hd__xnor2_1
  U767
  (
    .A(n870),
    .B(n795),
    .Y(n279)
  );


  sky130_fd_sc_hd__xor2_1
  U768
  (
    .A(n802),
    .B(n871),
    .X(n795)
  );


  sky130_fd_sc_hd__xor2_1
  U769
  (
    .A(n872),
    .B(n852),
    .X(n871)
  );


  sky130_fd_sc_hd__nor2_1
  U770
  (
    .A(n873),
    .B(n739),
    .Y(n852)
  );


  sky130_fd_sc_hd__xnor2_1
  U771
  (
    .A(n857),
    .B(n858),
    .Y(n870)
  );


  sky130_fd_sc_hd__xnor2_1
  U772
  (
    .A(n739),
    .B(n803),
    .Y(n858)
  );


  sky130_fd_sc_hd__a221oi_1
  U773
  (
    .A1(n783),
    .A2(n807),
    .B1(n874),
    .B2(n771),
    .C1(n875),
    .Y(n803)
  );


  sky130_fd_sc_hd__o22ai_1
  U774
  (
    .A1(n876),
    .A2(n787),
    .B1(n815),
    .B2(n789),
    .Y(n875)
  );


  sky130_fd_sc_hd__o22a_1
  U775
  (
    .A1(n801),
    .A2(n800),
    .B1(n802),
    .B2(n877),
    .X(n857)
  );


  sky130_fd_sc_hd__nor2_1
  U776
  (
    .A(n798),
    .B(n797),
    .Y(n877)
  );


  sky130_fd_sc_hd__xnor2_1
  U777
  (
    .A(n276),
    .B(n277),
    .Y(n869)
  );


  sky130_fd_sc_hd__xnor2_1
  U778
  (
    .A(n751),
    .B(n825),
    .Y(n277)
  );


  sky130_fd_sc_hd__a221oi_1
  U779
  (
    .A1(n878),
    .A2(n741),
    .B1(n862),
    .B2(n784),
    .C1(n879),
    .Y(n825)
  );


  sky130_fd_sc_hd__o22ai_1
  U780
  (
    .A1(n786),
    .A2(n811),
    .B1(n788),
    .B2(n880),
    .Y(n879)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U781
  (
    .B1(n881),
    .B2(n882),
    .A1_N(n883),
    .A2_N(n827),
    .Y(n276)
  );


  sky130_fd_sc_hd__nor2_1
  U782
  (
    .A(n881),
    .B(n882),
    .Y(n883)
  );


  sky130_fd_sc_hd__maj3_1
  U783
  (
    .A(n884),
    .B(n51),
    .C(n885),
    .X(n863)
  );


  sky130_fd_sc_hd__maj3_1
  U784
  (
    .A(n886),
    .B(n271),
    .C(n887),
    .X(n885)
  );


  sky130_fd_sc_hd__maj3_1
  U785
  (
    .A(n888),
    .B(n889),
    .C(n890),
    .X(n887)
  );


  sky130_fd_sc_hd__xor2_1
  U786
  (
    .A(n780),
    .B(n891),
    .X(n890)
  );


  sky130_fd_sc_hd__maj3_1
  U787
  (
    .A(n892),
    .B(n893),
    .C(n894),
    .X(n888)
  );


  sky130_fd_sc_hd__xor2_1
  U788
  (
    .A(n740),
    .B(n895),
    .X(n894)
  );


  sky130_fd_sc_hd__xor2_1
  U789
  (
    .A(n780),
    .B(n896),
    .X(n892)
  );


  sky130_fd_sc_hd__xor2_1
  U790
  (
    .A(n872),
    .B(n897),
    .X(n886)
  );


  sky130_fd_sc_hd__xnor2_1
  U791
  (
    .A(n898),
    .B(n272),
    .Y(n51)
  );


  sky130_fd_sc_hd__xor2_1
  U792
  (
    .A(n751),
    .B(n868),
    .X(n272)
  );


  sky130_fd_sc_hd__a221oi_1
  U793
  (
    .A1(n806),
    .A2(n862),
    .B1(n860),
    .B2(n807),
    .C1(n899),
    .Y(n868)
  );


  sky130_fd_sc_hd__o22ai_1
  U794
  (
    .A1(n786),
    .A2(n880),
    .B1(n788),
    .B2(n900),
    .Y(n899)
  );


  sky130_fd_sc_hd__xnor2_1
  U795
  (
    .A(n275),
    .B(n273),
    .Y(n898)
  );


  sky130_fd_sc_hd__xnor2_1
  U796
  (
    .A(n867),
    .B(n851),
    .Y(n273)
  );


  sky130_fd_sc_hd__o22ai_1
  U797
  (
    .A1(n901),
    .A2(n810),
    .B1(n902),
    .B2(n813),
    .Y(n867)
  );


  sky130_fd_sc_hd__xnor2_1
  U798
  (
    .A(n903),
    .B(n827),
    .Y(n275)
  );


  sky130_fd_sc_hd__xnor2_1
  U799
  (
    .A(n800),
    .B(n904),
    .Y(n827)
  );


  sky130_fd_sc_hd__xor2_1
  U800
  (
    .A(n798),
    .B(n802),
    .X(n904)
  );


  sky130_fd_sc_hd__clkinv_1
  U801
  (
    .A(n801),
    .Y(n798)
  );


  sky130_fd_sc_hd__nand2_1
  U802
  (
    .A(n740),
    .B(n905),
    .Y(n801)
  );


  sky130_fd_sc_hd__clkinv_1
  U803
  (
    .A(n797),
    .Y(n800)
  );


  sky130_fd_sc_hd__xor2_1
  U804
  (
    .A(n739),
    .B(n906),
    .X(n797)
  );


  sky130_fd_sc_hd__a221oi_1
  U805
  (
    .A1(n907),
    .A2(n771),
    .B1(n767),
    .B2(n908),
    .C1(n909),
    .Y(n906)
  );


  sky130_fd_sc_hd__o22ai_1
  U806
  (
    .A1(n876),
    .A2(n789),
    .B1(n815),
    .B2(n809),
    .Y(n909)
  );


  sky130_fd_sc_hd__xnor2_1
  U807
  (
    .A(n882),
    .B(n881),
    .Y(n903)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U808
  (
    .B1(n802),
    .B2(n910),
    .A1_N(n911),
    .A2_N(n912),
    .Y(n881)
  );


  sky130_fd_sc_hd__nor2_1
  U809
  (
    .A(n912),
    .B(n911),
    .Y(n910)
  );


  sky130_fd_sc_hd__o22ai_1
  U810
  (
    .A1(n913),
    .A2(n914),
    .B1(n915),
    .B2(n837),
    .Y(n882)
  );


  sky130_fd_sc_hd__and2_0
  U811
  (
    .A(n914),
    .B(n913),
    .X(n915)
  );


  sky130_fd_sc_hd__maj3_1
  U812
  (
    .A(n916),
    .B(n40),
    .C(n917),
    .X(n884)
  );


  sky130_fd_sc_hd__maj3_1
  U813
  (
    .A(n918),
    .B(n267),
    .C(n919),
    .X(n917)
  );


  sky130_fd_sc_hd__xor2_1
  U814
  (
    .A(n872),
    .B(n920),
    .X(n919)
  );


  sky130_fd_sc_hd__maj3_1
  U815
  (
    .A(n921),
    .B(n922),
    .C(n923),
    .X(n918)
  );


  sky130_fd_sc_hd__maj3_1
  U816
  (
    .A(n924),
    .B(n925),
    .C(n926),
    .X(n923)
  );


  sky130_fd_sc_hd__maj3_1
  U817
  (
    .A(n927),
    .B(n928),
    .C(n929),
    .X(n926)
  );


  sky130_fd_sc_hd__xor2_1
  U818
  (
    .A(n740),
    .B(n930),
    .X(n929)
  );


  sky130_fd_sc_hd__a21oi_1
  U819
  (
    .A1(n931),
    .A2(n932),
    .B1(n933),
    .Y(n927)
  );


  sky130_fd_sc_hd__o21a_1
  U820
  (
    .A1(n932),
    .A2(n931),
    .B1(A[15]),
    .X(n933)
  );


  sky130_fd_sc_hd__xor2_1
  U821
  (
    .A(n780),
    .B(n934),
    .X(n924)
  );


  sky130_fd_sc_hd__maj3_1
  U822
  (
    .A(n935),
    .B(n936),
    .C(n937),
    .X(n921)
  );


  sky130_fd_sc_hd__maj3_1
  U823
  (
    .A(n938),
    .B(n939),
    .C(n940),
    .X(n937)
  );


  sky130_fd_sc_hd__xor2_1
  U824
  (
    .A(n780),
    .B(n941),
    .X(n940)
  );


  sky130_fd_sc_hd__maj3_1
  U825
  (
    .A(n942),
    .B(n943),
    .C(n944),
    .X(n938)
  );


  sky130_fd_sc_hd__a21oi_1
  U826
  (
    .A1(n945),
    .A2(n946),
    .B1(n947),
    .Y(n944)
  );


  sky130_fd_sc_hd__a21oi_1
  U827
  (
    .A1(n948),
    .A2(n949),
    .B1(n97),
    .Y(n947)
  );


  sky130_fd_sc_hd__maj3_1
  U828
  (
    .A(n950),
    .B(n951),
    .C(n952),
    .X(n942)
  );


  sky130_fd_sc_hd__a21oi_1
  U829
  (
    .A1(n953),
    .A2(n954),
    .B1(n955),
    .Y(n952)
  );


  sky130_fd_sc_hd__a21oi_1
  U830
  (
    .A1(n956),
    .A2(n957),
    .B1(n97),
    .Y(n955)
  );


  sky130_fd_sc_hd__maj3_1
  U831
  (
    .A(n958),
    .B(n959),
    .C(n960),
    .X(n950)
  );


  sky130_fd_sc_hd__xor2_1
  U832
  (
    .A(n780),
    .B(n961),
    .X(n960)
  );


  sky130_fd_sc_hd__maj3_1
  U833
  (
    .A(n962),
    .B(n963),
    .C(n964),
    .X(n958)
  );


  sky130_fd_sc_hd__xor2_1
  U834
  (
    .A(n740),
    .B(n965),
    .X(n964)
  );


  sky130_fd_sc_hd__xor2_1
  U835
  (
    .A(n872),
    .B(n966),
    .X(n935)
  );


  sky130_fd_sc_hd__xnor2_1
  U836
  (
    .A(n967),
    .B(n271),
    .Y(n40)
  );


  sky130_fd_sc_hd__xnor2_1
  U837
  (
    .A(n968),
    .B(n837),
    .Y(n271)
  );


  sky130_fd_sc_hd__xnor2_1
  U838
  (
    .A(n912),
    .B(n969),
    .Y(n837)
  );


  sky130_fd_sc_hd__xnor2_1
  U839
  (
    .A(n802),
    .B(n911),
    .Y(n969)
  );


  sky130_fd_sc_hd__maj3_1
  U840
  (
    .A(n832),
    .B(n834),
    .C(n831),
    .X(n911)
  );


  sky130_fd_sc_hd__nor2_1
  U841
  (
    .A(n970),
    .B(n739),
    .Y(n802)
  );


  sky130_fd_sc_hd__xnor2_1
  U842
  (
    .A(n740),
    .B(n835),
    .Y(n912)
  );


  sky130_fd_sc_hd__a221oi_1
  U843
  (
    .A1(n971),
    .A2(n771),
    .B1(n767),
    .B2(n905),
    .C1(n972),
    .Y(n835)
  );


  sky130_fd_sc_hd__o22ai_1
  U844
  (
    .A1(n873),
    .A2(n789),
    .B1(n876),
    .B2(n809),
    .Y(n972)
  );


  sky130_fd_sc_hd__xnor2_1
  U845
  (
    .A(n914),
    .B(n913),
    .Y(n968)
  );


  sky130_fd_sc_hd__o22a_1
  U846
  (
    .A1(n973),
    .A2(n974),
    .B1(n975),
    .B2(n840),
    .X(n913)
  );


  sky130_fd_sc_hd__and2_0
  U847
  (
    .A(n974),
    .B(n973),
    .X(n975)
  );


  sky130_fd_sc_hd__xnor2_1
  U848
  (
    .A(n751),
    .B(n848),
    .Y(n914)
  );


  sky130_fd_sc_hd__a221oi_1
  U849
  (
    .A1(n861),
    .A2(n807),
    .B1(n855),
    .B2(n862),
    .C1(n976),
    .Y(n848)
  );


  sky130_fd_sc_hd__o22ai_1
  U850
  (
    .A1(n815),
    .A2(n811),
    .B1(n786),
    .B2(n900),
    .Y(n976)
  );


  sky130_fd_sc_hd__xnor2_1
  U851
  (
    .A(n269),
    .B(n268),
    .Y(n967)
  );


  sky130_fd_sc_hd__o22a_1
  U852
  (
    .A1(n977),
    .A2(n978),
    .B1(n979),
    .B2(n889),
    .X(n268)
  );


  sky130_fd_sc_hd__and2_0
  U853
  (
    .A(n978),
    .B(n977),
    .X(n979)
  );


  sky130_fd_sc_hd__xnor2_1
  U854
  (
    .A(n851),
    .B(n897),
    .Y(n269)
  );


  sky130_fd_sc_hd__a222oi_1
  U855
  (
    .A1(n980),
    .A2(n768),
    .B1(n741),
    .B2(n981),
    .C1(n770),
    .C2(n982),
    .Y(n897)
  );


  sky130_fd_sc_hd__maj3_1
  U856
  (
    .A(n983),
    .B(n30),
    .C(n984),
    .X(n916)
  );


  sky130_fd_sc_hd__maj3_1
  U857
  (
    .A(n985),
    .B(n263),
    .C(n986),
    .X(n984)
  );


  sky130_fd_sc_hd__xor2_1
  U858
  (
    .A(n834),
    .B(n987),
    .X(n986)
  );


  sky130_fd_sc_hd__xor2_1
  U859
  (
    .A(n872),
    .B(n988),
    .X(n985)
  );


  sky130_fd_sc_hd__xnor2_1
  U860
  (
    .A(n989),
    .B(n267),
    .Y(n30)
  );


  sky130_fd_sc_hd__xnor2_1
  U861
  (
    .A(n990),
    .B(n889),
    .Y(n267)
  );


  sky130_fd_sc_hd__xnor2_1
  U862
  (
    .A(n991),
    .B(n840),
    .Y(n889)
  );


  sky130_fd_sc_hd__xor2_1
  U863
  (
    .A(n832),
    .B(n992),
    .X(n840)
  );


  sky130_fd_sc_hd__xor2_1
  U864
  (
    .A(A[9]),
    .B(n831),
    .X(n992)
  );


  sky130_fd_sc_hd__nor2_1
  U865
  (
    .A(n993),
    .B(n739),
    .Y(n831)
  );


  sky130_fd_sc_hd__xnor2_1
  U866
  (
    .A(n974),
    .B(n973),
    .Y(n991)
  );


  sky130_fd_sc_hd__o22a_1
  U867
  (
    .A1(n846),
    .A2(n847),
    .B1(n832),
    .B2(n994),
    .X(n973)
  );


  sky130_fd_sc_hd__nor2_1
  U868
  (
    .A(n843),
    .B(n844),
    .Y(n994)
  );


  sky130_fd_sc_hd__xnor2_1
  U869
  (
    .A(n739),
    .B(n842),
    .Y(n974)
  );


  sky130_fd_sc_hd__a221oi_1
  U870
  (
    .A1(n769),
    .A2(n905),
    .B1(n995),
    .B2(n771),
    .C1(n996),
    .Y(n842)
  );


  sky130_fd_sc_hd__o22ai_1
  U871
  (
    .A1(n970),
    .A2(n787),
    .B1(n873),
    .B2(n809),
    .Y(n996)
  );


  sky130_fd_sc_hd__xnor2_1
  U872
  (
    .A(n977),
    .B(n978),
    .Y(n990)
  );


  sky130_fd_sc_hd__xnor2_1
  U873
  (
    .A(n751),
    .B(n891),
    .Y(n978)
  );


  sky130_fd_sc_hd__a221oi_1
  U874
  (
    .A1(n878),
    .A2(n807),
    .B1(n874),
    .B2(n862),
    .C1(n997),
    .Y(n891)
  );


  sky130_fd_sc_hd__o22ai_1
  U875
  (
    .A1(n876),
    .A2(n811),
    .B1(n815),
    .B2(n880),
    .Y(n997)
  );


  sky130_fd_sc_hd__o22a_1
  U876
  (
    .A1(n998),
    .A2(n999),
    .B1(n1000),
    .B2(n893),
    .X(n977)
  );


  sky130_fd_sc_hd__and2_0
  U877
  (
    .A(n999),
    .B(n998),
    .X(n1000)
  );


  sky130_fd_sc_hd__xnor2_1
  U878
  (
    .A(n264),
    .B(n265),
    .Y(n989)
  );


  sky130_fd_sc_hd__xnor2_1
  U879
  (
    .A(n851),
    .B(n920),
    .Y(n265)
  );


  sky130_fd_sc_hd__a221oi_1
  U880
  (
    .A1(n741),
    .A2(n1001),
    .B1(n982),
    .B2(n784),
    .C1(n1002),
    .Y(n920)
  );


  sky130_fd_sc_hd__o22ai_1
  U881
  (
    .A1(n901),
    .A2(n786),
    .B1(n1003),
    .B2(n788),
    .Y(n1002)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U882
  (
    .B1(n1004),
    .B2(n1005),
    .A1_N(n1006),
    .A2_N(n922),
    .Y(n264)
  );


  sky130_fd_sc_hd__nor2_1
  U883
  (
    .A(n1005),
    .B(n1004),
    .Y(n1006)
  );


  sky130_fd_sc_hd__maj3_1
  U884
  (
    .A(n1007),
    .B(n257),
    .C(n1008),
    .X(n983)
  );


  sky130_fd_sc_hd__maj3_1
  U885
  (
    .A(n1009),
    .B(n395),
    .C(n1010),
    .X(n1008)
  );


  sky130_fd_sc_hd__maj3_1
  U886
  (
    .A(n1011),
    .B(n1012),
    .C(n1013),
    .X(n1010)
  );


  sky130_fd_sc_hd__xor2_1
  U887
  (
    .A(n872),
    .B(n1014),
    .X(n1013)
  );


  sky130_fd_sc_hd__maj3_1
  U888
  (
    .A(n1015),
    .B(n1016),
    .C(n1017),
    .X(n1011)
  );


  sky130_fd_sc_hd__xor2_1
  U889
  (
    .A(n780),
    .B(n1018),
    .X(n1017)
  );


  sky130_fd_sc_hd__xor2_1
  U890
  (
    .A(n872),
    .B(n1019),
    .X(n1015)
  );


  sky130_fd_sc_hd__xor2_1
  U891
  (
    .A(A[9]),
    .B(n1020),
    .X(n1009)
  );


  sky130_fd_sc_hd__xnor2_1
  U892
  (
    .A(n1021),
    .B(n261),
    .Y(n257)
  );


  sky130_fd_sc_hd__xor2_1
  U893
  (
    .A(n987),
    .B(A[9]),
    .X(n261)
  );


  sky130_fd_sc_hd__o22ai_1
  U894
  (
    .A1(n810),
    .A2(n1022),
    .B1(n1023),
    .B2(n813),
    .Y(n987)
  );


  sky130_fd_sc_hd__xnor2_1
  U895
  (
    .A(n263),
    .B(n260),
    .Y(n1021)
  );


  sky130_fd_sc_hd__xnor2_1
  U896
  (
    .A(n872),
    .B(n988),
    .Y(n260)
  );


  sky130_fd_sc_hd__a221oi_1
  U897
  (
    .A1(n806),
    .A2(n982),
    .B1(n807),
    .B2(n980),
    .C1(n1024),
    .Y(n988)
  );


  sky130_fd_sc_hd__o22ai_1
  U898
  (
    .A1(n1003),
    .A2(n786),
    .B1(n788),
    .B2(n1025),
    .Y(n1024)
  );


  sky130_fd_sc_hd__xnor2_1
  U899
  (
    .A(n1026),
    .B(n922),
    .Y(n263)
  );


  sky130_fd_sc_hd__xnor2_1
  U900
  (
    .A(n1027),
    .B(n893),
    .Y(n922)
  );


  sky130_fd_sc_hd__xnor2_1
  U901
  (
    .A(n846),
    .B(n1028),
    .Y(n893)
  );


  sky130_fd_sc_hd__xor2_1
  U902
  (
    .A(n832),
    .B(n843),
    .X(n1028)
  );


  sky130_fd_sc_hd__nor2_1
  U903
  (
    .A(n1029),
    .B(n739),
    .Y(n832)
  );


  sky130_fd_sc_hd__clkinv_1
  U904
  (
    .A(n844),
    .Y(n846)
  );


  sky130_fd_sc_hd__o22ai_1
  U905
  (
    .A1(n1030),
    .A2(n1031),
    .B1(n843),
    .B2(n1032),
    .Y(n844)
  );


  sky130_fd_sc_hd__nor2_1
  U906
  (
    .A(n1033),
    .B(n1034),
    .Y(n1032)
  );


  sky130_fd_sc_hd__xnor2_1
  U907
  (
    .A(n998),
    .B(n999),
    .Y(n1027)
  );


  sky130_fd_sc_hd__xnor2_1
  U908
  (
    .A(n739),
    .B(n895),
    .Y(n999)
  );


  sky130_fd_sc_hd__a221oi_1
  U909
  (
    .A1(n1035),
    .A2(n771),
    .B1(n767),
    .B2(B[9]),
    .C1(n1036),
    .Y(n895)
  );


  sky130_fd_sc_hd__o22ai_1
  U910
  (
    .A1(n970),
    .A2(n789),
    .B1(n1037),
    .B2(n809),
    .Y(n1036)
  );


  sky130_fd_sc_hd__xnor2_1
  U911
  (
    .A(n751),
    .B(n896),
    .Y(n998)
  );


  sky130_fd_sc_hd__a221oi_1
  U912
  (
    .A1(n907),
    .A2(n862),
    .B1(n860),
    .B2(n908),
    .C1(n1038),
    .Y(n896)
  );


  sky130_fd_sc_hd__o22ai_1
  U913
  (
    .A1(n876),
    .A2(n880),
    .B1(n815),
    .B2(n900),
    .Y(n1038)
  );


  sky130_fd_sc_hd__xnor2_1
  U914
  (
    .A(n1005),
    .B(n1004),
    .Y(n1026)
  );


  sky130_fd_sc_hd__o22ai_1
  U915
  (
    .A1(n1039),
    .A2(n1040),
    .B1(n1041),
    .B2(n925),
    .Y(n1004)
  );


  sky130_fd_sc_hd__nor2_1
  U916
  (
    .A(n1042),
    .B(n1043),
    .Y(n1041)
  );


  sky130_fd_sc_hd__clkinv_1
  U917
  (
    .A(n1042),
    .Y(n1040)
  );


  sky130_fd_sc_hd__o22ai_1
  U918
  (
    .A1(n1044),
    .A2(n1045),
    .B1(n1046),
    .B2(n936),
    .Y(n1005)
  );


  sky130_fd_sc_hd__nor2_1
  U919
  (
    .A(n1047),
    .B(n1048),
    .Y(n1046)
  );


  sky130_fd_sc_hd__clkinv_1
  U920
  (
    .A(n1047),
    .Y(n1045)
  );


  sky130_fd_sc_hd__maj3_1
  U921
  (
    .A(n1049),
    .B(n362),
    .C(n1050),
    .X(n1007)
  );


  sky130_fd_sc_hd__maj3_1
  U922
  (
    .A(n1051),
    .B(n402),
    .C(n1052),
    .X(n1050)
  );


  sky130_fd_sc_hd__xor2_1
  U923
  (
    .A(A[9]),
    .B(n1053),
    .X(n1052)
  );


  sky130_fd_sc_hd__maj3_1
  U924
  (
    .A(n1054),
    .B(n1055),
    .C(n1056),
    .X(n1051)
  );


  sky130_fd_sc_hd__maj3_1
  U925
  (
    .A(n1057),
    .B(n1058),
    .C(n1059),
    .X(n1056)
  );


  sky130_fd_sc_hd__xor2_1
  U926
  (
    .A(n780),
    .B(n1060),
    .X(n1059)
  );


  sky130_fd_sc_hd__xor2_1
  U927
  (
    .A(n872),
    .B(n1061),
    .X(n1057)
  );


  sky130_fd_sc_hd__maj3_1
  U928
  (
    .A(n1062),
    .B(n1063),
    .C(n1064),
    .X(n1054)
  );


  sky130_fd_sc_hd__maj3_1
  U929
  (
    .A(n1065),
    .B(n1066),
    .C(n1067),
    .X(n1064)
  );


  sky130_fd_sc_hd__xor2_1
  U930
  (
    .A(n872),
    .B(n1068),
    .X(n1067)
  );


  sky130_fd_sc_hd__maj3_1
  U931
  (
    .A(n1069),
    .B(n1070),
    .C(n1071),
    .X(n1065)
  );


  sky130_fd_sc_hd__xor2_1
  U932
  (
    .A(n780),
    .B(n1072),
    .X(n1071)
  );


  sky130_fd_sc_hd__maj3_1
  U933
  (
    .A(n1073),
    .B(n1074),
    .C(n1075),
    .X(n1069)
  );


  sky130_fd_sc_hd__xor2_1
  U934
  (
    .A(n780),
    .B(n1076),
    .X(n1075)
  );


  sky130_fd_sc_hd__maj3_1
  U935
  (
    .A(n1077),
    .B(n1078),
    .C(n1079),
    .X(n1073)
  );


  sky130_fd_sc_hd__xor2_1
  U936
  (
    .A(n780),
    .B(n1080),
    .X(n1079)
  );


  sky130_fd_sc_hd__maj3_1
  U937
  (
    .A(n1081),
    .B(n1082),
    .C(n1083),
    .X(n1077)
  );


  sky130_fd_sc_hd__xor2_1
  U938
  (
    .A(n780),
    .B(n1084),
    .X(n1083)
  );


  sky130_fd_sc_hd__maj3_1
  U939
  (
    .A(n1085),
    .B(n1086),
    .C(n1087),
    .X(n1062)
  );


  sky130_fd_sc_hd__xor2_1
  U940
  (
    .A(A[9]),
    .B(n1088),
    .X(n1087)
  );


  sky130_fd_sc_hd__maj3_1
  U941
  (
    .A(n1089),
    .B(n1090),
    .C(n1091),
    .X(n1085)
  );


  sky130_fd_sc_hd__xor2_1
  U942
  (
    .A(n872),
    .B(n1092),
    .X(n1091)
  );


  sky130_fd_sc_hd__maj3_1
  U943
  (
    .A(n1093),
    .B(n1094),
    .C(n1095),
    .X(n1089)
  );


  sky130_fd_sc_hd__xor2_1
  U944
  (
    .A(n872),
    .B(n1096),
    .X(n1095)
  );


  sky130_fd_sc_hd__maj3_1
  U945
  (
    .A(n1097),
    .B(n1098),
    .C(n1099),
    .X(n1093)
  );


  sky130_fd_sc_hd__xor2_1
  U946
  (
    .A(n872),
    .B(n1100),
    .X(n1099)
  );


  sky130_fd_sc_hd__maj3_1
  U947
  (
    .A(n1101),
    .B(n1102),
    .C(n1103),
    .X(n1097)
  );


  sky130_fd_sc_hd__xor2_1
  U948
  (
    .A(n872),
    .B(n1104),
    .X(n1103)
  );


  sky130_fd_sc_hd__maj3_1
  U949
  (
    .A(n1105),
    .B(n1106),
    .C(n1107),
    .X(n1101)
  );


  sky130_fd_sc_hd__xor2_1
  U950
  (
    .A(n872),
    .B(n1108),
    .X(n1107)
  );


  sky130_fd_sc_hd__maj3_1
  U951
  (
    .A(n1109),
    .B(n1110),
    .C(n1111),
    .X(n1105)
  );


  sky130_fd_sc_hd__xor2_1
  U952
  (
    .A(n872),
    .B(n1112),
    .X(n1111)
  );


  sky130_fd_sc_hd__maj3_1
  U953
  (
    .A(n1113),
    .B(n1114),
    .C(n1115),
    .X(n1109)
  );


  sky130_fd_sc_hd__xor2_1
  U954
  (
    .A(n872),
    .B(n1116),
    .X(n1115)
  );


  sky130_fd_sc_hd__xnor2_1
  U955
  (
    .A(n1117),
    .B(n395),
    .Y(n362)
  );


  sky130_fd_sc_hd__xnor2_1
  U956
  (
    .A(n1118),
    .B(n936),
    .Y(n395)
  );


  sky130_fd_sc_hd__xnor2_1
  U957
  (
    .A(n1119),
    .B(n925),
    .Y(n936)
  );


  sky130_fd_sc_hd__xor2_1
  U958
  (
    .A(n1031),
    .B(n1120),
    .X(n925)
  );


  sky130_fd_sc_hd__xor2_1
  U959
  (
    .A(n843),
    .B(n1030),
    .X(n1120)
  );


  sky130_fd_sc_hd__clkinv_1
  U960
  (
    .A(n1034),
    .Y(n1030)
  );


  sky130_fd_sc_hd__o22ai_1
  U961
  (
    .A1(A[12]),
    .A2(n1121),
    .B1(A[15]),
    .B2(n1122),
    .Y(n1034)
  );


  sky130_fd_sc_hd__and2_0
  U962
  (
    .A(n1121),
    .B(A[12]),
    .X(n1122)
  );


  sky130_fd_sc_hd__clkinv_1
  U963
  (
    .A(n847),
    .Y(n843)
  );


  sky130_fd_sc_hd__nand2_1
  U964
  (
    .A(n740),
    .B(B[11]),
    .Y(n847)
  );


  sky130_fd_sc_hd__clkinv_1
  U965
  (
    .A(n1033),
    .Y(n1031)
  );


  sky130_fd_sc_hd__xor2_1
  U966
  (
    .A(n739),
    .B(n1123),
    .X(n1033)
  );


  sky130_fd_sc_hd__a221oi_1
  U967
  (
    .A1(n769),
    .A2(B[9]),
    .B1(n1124),
    .B2(n771),
    .C1(n1125),
    .Y(n1123)
  );


  sky130_fd_sc_hd__o22ai_1
  U968
  (
    .A1(n1029),
    .A2(n787),
    .B1(n970),
    .B2(n809),
    .Y(n1125)
  );


  sky130_fd_sc_hd__xor2_1
  U969
  (
    .A(n1042),
    .B(n1039),
    .X(n1119)
  );


  sky130_fd_sc_hd__clkinv_1
  U970
  (
    .A(n1043),
    .Y(n1039)
  );


  sky130_fd_sc_hd__o22ai_1
  U971
  (
    .A1(n1126),
    .A2(n1127),
    .B1(n1128),
    .B2(n928),
    .Y(n1043)
  );


  sky130_fd_sc_hd__and2_0
  U972
  (
    .A(n1127),
    .B(n1126),
    .X(n1128)
  );


  sky130_fd_sc_hd__xor2_1
  U973
  (
    .A(n751),
    .B(n934),
    .X(n1042)
  );


  sky130_fd_sc_hd__a221oi_1
  U974
  (
    .A1(n862),
    .A2(n971),
    .B1(n860),
    .B2(n905),
    .C1(n1129),
    .Y(n934)
  );


  sky130_fd_sc_hd__o22ai_1
  U975
  (
    .A1(n873),
    .A2(n880),
    .B1(n876),
    .B2(n900),
    .Y(n1129)
  );


  sky130_fd_sc_hd__xor2_1
  U976
  (
    .A(n1047),
    .B(n1044),
    .X(n1118)
  );


  sky130_fd_sc_hd__clkinv_1
  U977
  (
    .A(n1048),
    .Y(n1044)
  );


  sky130_fd_sc_hd__o22ai_1
  U978
  (
    .A1(n1130),
    .A2(n1131),
    .B1(n1132),
    .B2(n939),
    .Y(n1048)
  );


  sky130_fd_sc_hd__and2_0
  U979
  (
    .A(n1131),
    .B(n1130),
    .X(n1132)
  );


  sky130_fd_sc_hd__xor2_1
  U980
  (
    .A(n851),
    .B(n966),
    .X(n1047)
  );


  sky130_fd_sc_hd__a221oi_1
  U981
  (
    .A1(n807),
    .A2(n981),
    .B1(n855),
    .B2(n982),
    .C1(n1133),
    .Y(n966)
  );


  sky130_fd_sc_hd__o22ai_1
  U982
  (
    .A1(n901),
    .A2(n815),
    .B1(n786),
    .B2(n1025),
    .Y(n1133)
  );


  sky130_fd_sc_hd__xor2_1
  U983
  (
    .A(n396),
    .B(n392),
    .X(n1117)
  );


  sky130_fd_sc_hd__clkinv_1
  U984
  (
    .A(n397),
    .Y(n392)
  );


  sky130_fd_sc_hd__o22ai_1
  U985
  (
    .A1(n1134),
    .A2(n1135),
    .B1(n1136),
    .B2(n1012),
    .Y(n397)
  );


  sky130_fd_sc_hd__and2_0
  U986
  (
    .A(n1135),
    .B(n1134),
    .X(n1136)
  );


  sky130_fd_sc_hd__xor2_1
  U987
  (
    .A(n834),
    .B(n1020),
    .X(n396)
  );


  sky130_fd_sc_hd__a222oi_1
  U988
  (
    .A1(n1137),
    .A2(n768),
    .B1(n1138),
    .B2(n741),
    .C1(n770),
    .C2(n1139),
    .Y(n1020)
  );


  sky130_fd_sc_hd__maj3_1
  U989
  (
    .A(n1140),
    .B(n349),
    .C(n1141),
    .X(n1049)
  );


  sky130_fd_sc_hd__maj3_1
  U990
  (
    .A(n1142),
    .B(n458),
    .C(n1143),
    .X(n1141)
  );


  sky130_fd_sc_hd__xor2_1
  U991
  (
    .A(A[9]),
    .B(n1144),
    .X(n1143)
  );


  sky130_fd_sc_hd__xor2_1
  U992
  (
    .A(n1145),
    .B(n1146),
    .X(n1142)
  );


  sky130_fd_sc_hd__xnor2_1
  U993
  (
    .A(n1147),
    .B(n402),
    .Y(n349)
  );


  sky130_fd_sc_hd__xnor2_1
  U994
  (
    .A(n1148),
    .B(n1012),
    .Y(n402)
  );


  sky130_fd_sc_hd__xnor2_1
  U995
  (
    .A(n1149),
    .B(n939),
    .Y(n1012)
  );


  sky130_fd_sc_hd__xnor2_1
  U996
  (
    .A(n1150),
    .B(n928),
    .Y(n939)
  );


  sky130_fd_sc_hd__xnor2_1
  U997
  (
    .A(n1151),
    .B(n1121),
    .Y(n928)
  );


  sky130_fd_sc_hd__nand2_1
  U998
  (
    .A(n740),
    .B(B[12]),
    .Y(n1121)
  );


  sky130_fd_sc_hd__xor2_1
  U999
  (
    .A(n1145),
    .B(A[15]),
    .X(n1151)
  );


  sky130_fd_sc_hd__xnor2_1
  U1000
  (
    .A(n1126),
    .B(n1127),
    .Y(n1150)
  );


  sky130_fd_sc_hd__xnor2_1
  U1001
  (
    .A(n739),
    .B(n930),
    .Y(n1127)
  );


  sky130_fd_sc_hd__a221oi_1
  U1002
  (
    .A1(n783),
    .A2(B[9]),
    .B1(n1152),
    .B2(n771),
    .C1(n1153),
    .Y(n930)
  );


  sky130_fd_sc_hd__o22ai_1
  U1003
  (
    .A1(n1154),
    .A2(n787),
    .B1(n1029),
    .B2(n789),
    .Y(n1153)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1004
  (
    .B1(n932),
    .B2(n931),
    .A1_N(n1155),
    .A2_N(n97),
    .Y(n1126)
  );


  sky130_fd_sc_hd__nor2_1
  U1005
  (
    .A(n931),
    .B(n932),
    .Y(n1155)
  );


  sky130_fd_sc_hd__xnor2_1
  U1006
  (
    .A(n1130),
    .B(n1131),
    .Y(n1149)
  );


  sky130_fd_sc_hd__xnor2_1
  U1007
  (
    .A(n751),
    .B(n941),
    .Y(n1131)
  );


  sky130_fd_sc_hd__a221oi_1
  U1008
  (
    .A1(n861),
    .A2(n905),
    .B1(n995),
    .B2(n862),
    .C1(n1156),
    .Y(n941)
  );


  sky130_fd_sc_hd__o22ai_1
  U1009
  (
    .A1(n970),
    .A2(n811),
    .B1(n873),
    .B2(n900),
    .Y(n1156)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1010
  (
    .B1(n1157),
    .B2(n1158),
    .A1_N(n1159),
    .A2_N(n943),
    .Y(n1130)
  );


  sky130_fd_sc_hd__nor2_1
  U1011
  (
    .A(n1158),
    .B(n1157),
    .Y(n1159)
  );


  sky130_fd_sc_hd__xnor2_1
  U1012
  (
    .A(n1134),
    .B(n1135),
    .Y(n1148)
  );


  sky130_fd_sc_hd__xnor2_1
  U1013
  (
    .A(n851),
    .B(n1014),
    .Y(n1135)
  );


  sky130_fd_sc_hd__a221oi_1
  U1014
  (
    .A1(n807),
    .A2(n1001),
    .B1(n874),
    .B2(n982),
    .C1(n1160),
    .Y(n1014)
  );


  sky130_fd_sc_hd__o22ai_1
  U1015
  (
    .A1(n901),
    .A2(n876),
    .B1(n1003),
    .B2(n815),
    .Y(n1160)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1016
  (
    .B1(n1161),
    .B2(n1162),
    .A1_N(n1163),
    .A2_N(n1016),
    .Y(n1134)
  );


  sky130_fd_sc_hd__nor2_1
  U1017
  (
    .A(n1162),
    .B(n1161),
    .Y(n1163)
  );


  sky130_fd_sc_hd__xnor2_1
  U1018
  (
    .A(n399),
    .B(n400),
    .Y(n1147)
  );


  sky130_fd_sc_hd__xnor2_1
  U1019
  (
    .A(n834),
    .B(n1053),
    .Y(n400)
  );


  sky130_fd_sc_hd__a221oi_1
  U1020
  (
    .A1(n1164),
    .A2(n741),
    .B1(n1139),
    .B2(n784),
    .C1(n1165),
    .Y(n1053)
  );


  sky130_fd_sc_hd__o22ai_1
  U1021
  (
    .A1(n786),
    .A2(n1022),
    .B1(n788),
    .B2(n1166),
    .Y(n1165)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1022
  (
    .B1(n1167),
    .B2(n1168),
    .A1_N(n1169),
    .A2_N(n1055),
    .Y(n399)
  );


  sky130_fd_sc_hd__nor2_1
  U1023
  (
    .A(n1168),
    .B(n1167),
    .Y(n1169)
  );


  sky130_fd_sc_hd__maj3_1
  U1024
  (
    .A(n1170),
    .B(n338),
    .C(n1171),
    .X(n1140)
  );


  sky130_fd_sc_hd__maj3_1
  U1025
  (
    .A(n1172),
    .B(n410),
    .C(n1173),
    .X(n1171)
  );


  sky130_fd_sc_hd__xor2_1
  U1026
  (
    .A(A[9]),
    .B(n1174),
    .X(n1173)
  );


  sky130_fd_sc_hd__xor2_1
  U1027
  (
    .A(A[12]),
    .B(n1175),
    .X(n1172)
  );


  sky130_fd_sc_hd__xnor2_1
  U1028
  (
    .A(n1176),
    .B(n456),
    .Y(n338)
  );


  sky130_fd_sc_hd__xnor2_1
  U1029
  (
    .A(n834),
    .B(n1144),
    .Y(n456)
  );


  sky130_fd_sc_hd__a221oi_1
  U1030
  (
    .A1(n806),
    .A2(n1139),
    .B1(n1137),
    .B2(n807),
    .C1(n1177),
    .Y(n1144)
  );


  sky130_fd_sc_hd__o22ai_1
  U1031
  (
    .A1(n786),
    .A2(n1166),
    .B1(n788),
    .B2(n1178),
    .Y(n1177)
  );


  sky130_fd_sc_hd__xnor2_1
  U1032
  (
    .A(n458),
    .B(n455),
    .Y(n1176)
  );


  sky130_fd_sc_hd__xnor2_1
  U1033
  (
    .A(n1146),
    .B(A[12]),
    .Y(n455)
  );


  sky130_fd_sc_hd__o22ai_1
  U1034
  (
    .A1(n810),
    .A2(n1179),
    .B1(n813),
    .B2(n1180),
    .Y(n1146)
  );


  sky130_fd_sc_hd__xnor2_1
  U1035
  (
    .A(n1181),
    .B(n1055),
    .Y(n458)
  );


  sky130_fd_sc_hd__xnor2_1
  U1036
  (
    .A(n1162),
    .B(n1182),
    .Y(n1055)
  );


  sky130_fd_sc_hd__xnor2_1
  U1037
  (
    .A(n1161),
    .B(n1016),
    .Y(n1182)
  );


  sky130_fd_sc_hd__xnor2_1
  U1038
  (
    .A(n1183),
    .B(n943),
    .Y(n1016)
  );


  sky130_fd_sc_hd__xnor2_1
  U1039
  (
    .A(n932),
    .B(n1184),
    .Y(n943)
  );


  sky130_fd_sc_hd__xor2_1
  U1040
  (
    .A(A[15]),
    .B(n931),
    .X(n1184)
  );


  sky130_fd_sc_hd__nor2_1
  U1041
  (
    .A(n739),
    .B(n1185),
    .Y(n931)
  );


  sky130_fd_sc_hd__xnor2_1
  U1042
  (
    .A(n740),
    .B(n1186),
    .Y(n932)
  );


  sky130_fd_sc_hd__a221oi_1
  U1043
  (
    .A1(n771),
    .A2(n1187),
    .B1(n767),
    .B2(B[12]),
    .C1(n1188),
    .Y(n1186)
  );


  sky130_fd_sc_hd__o22ai_1
  U1044
  (
    .A1(n1029),
    .A2(n809),
    .B1(n1154),
    .B2(n789),
    .Y(n1188)
  );


  sky130_fd_sc_hd__xnor2_1
  U1045
  (
    .A(n1158),
    .B(n1157),
    .Y(n1183)
  );


  sky130_fd_sc_hd__o22ai_1
  U1046
  (
    .A1(n948),
    .A2(n949),
    .B1(n1189),
    .B2(n97),
    .Y(n1157)
  );


  sky130_fd_sc_hd__nor2_1
  U1047
  (
    .A(n945),
    .B(n946),
    .Y(n1189)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1048
  (
    .B1(n1190),
    .B2(n951),
    .A1_N(n1191),
    .A2_N(n1192),
    .Y(n1158)
  );


  sky130_fd_sc_hd__nor2_1
  U1049
  (
    .A(n1192),
    .B(n1191),
    .Y(n1190)
  );


  sky130_fd_sc_hd__xor2_1
  U1050
  (
    .A(n751),
    .B(n1018),
    .X(n1161)
  );


  sky130_fd_sc_hd__a221oi_1
  U1051
  (
    .A1(n1035),
    .A2(n862),
    .B1(n860),
    .B2(B[9]),
    .C1(n1193),
    .Y(n1018)
  );


  sky130_fd_sc_hd__o22ai_1
  U1052
  (
    .A1(n970),
    .A2(n880),
    .B1(n1037),
    .B2(n900),
    .Y(n1193)
  );


  sky130_fd_sc_hd__xor2_1
  U1053
  (
    .A(n851),
    .B(n1019),
    .X(n1162)
  );


  sky130_fd_sc_hd__a221oi_1
  U1054
  (
    .A1(n907),
    .A2(n982),
    .B1(n908),
    .B2(n980),
    .C1(n1194),
    .Y(n1019)
  );


  sky130_fd_sc_hd__o22ai_1
  U1055
  (
    .A1(n1003),
    .A2(n876),
    .B1(n1025),
    .B2(n815),
    .Y(n1194)
  );


  sky130_fd_sc_hd__xnor2_1
  U1056
  (
    .A(n1168),
    .B(n1167),
    .Y(n1181)
  );


  sky130_fd_sc_hd__o22ai_1
  U1057
  (
    .A1(n1195),
    .A2(n1196),
    .B1(n1197),
    .B2(n1058),
    .Y(n1167)
  );


  sky130_fd_sc_hd__and2_0
  U1058
  (
    .A(n1196),
    .B(n1195),
    .X(n1197)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1059
  (
    .B1(n1198),
    .B2(n1063),
    .A1_N(n1199),
    .A2_N(n1200),
    .Y(n1168)
  );


  sky130_fd_sc_hd__nor2_1
  U1060
  (
    .A(n1200),
    .B(n1199),
    .Y(n1198)
  );


  sky130_fd_sc_hd__maj3_1
  U1061
  (
    .A(n1201),
    .B(n328),
    .C(n1202),
    .X(n1170)
  );


  sky130_fd_sc_hd__maj3_1
  U1062
  (
    .A(n1203),
    .B(n454),
    .C(n1204),
    .X(n1202)
  );


  sky130_fd_sc_hd__xor2_1
  U1063
  (
    .A(A[12]),
    .B(n1205),
    .X(n1204)
  );


  sky130_fd_sc_hd__maj3_1
  U1064
  (
    .A(n1206),
    .B(n1207),
    .C(n1208),
    .X(n1203)
  );


  sky130_fd_sc_hd__xor2_1
  U1065
  (
    .A(A[9]),
    .B(n1209),
    .X(n1208)
  );


  sky130_fd_sc_hd__maj3_1
  U1066
  (
    .A(n1210),
    .B(n1211),
    .C(n1212),
    .X(n1206)
  );


  sky130_fd_sc_hd__xor2_1
  U1067
  (
    .A(A[9]),
    .B(n1213),
    .X(n1212)
  );


  sky130_fd_sc_hd__maj3_1
  U1068
  (
    .A(n1214),
    .B(n1215),
    .C(n1216),
    .X(n1210)
  );


  sky130_fd_sc_hd__xor2_1
  U1069
  (
    .A(A[9]),
    .B(n1217),
    .X(n1216)
  );


  sky130_fd_sc_hd__maj3_1
  U1070
  (
    .A(n1218),
    .B(n1219),
    .C(n1220),
    .X(n1214)
  );


  sky130_fd_sc_hd__xor2_1
  U1071
  (
    .A(A[9]),
    .B(n1221),
    .X(n1220)
  );


  sky130_fd_sc_hd__maj3_1
  U1072
  (
    .A(n1222),
    .B(n1223),
    .C(n1224),
    .X(n1218)
  );


  sky130_fd_sc_hd__xor2_1
  U1073
  (
    .A(A[9]),
    .B(n1225),
    .X(n1224)
  );


  sky130_fd_sc_hd__maj3_1
  U1074
  (
    .A(n1226),
    .B(n1227),
    .C(n1228),
    .X(n1222)
  );


  sky130_fd_sc_hd__xor2_1
  U1075
  (
    .A(A[9]),
    .B(n1229),
    .X(n1228)
  );


  sky130_fd_sc_hd__maj3_1
  U1076
  (
    .A(n1230),
    .B(n1231),
    .C(n1232),
    .X(n1226)
  );


  sky130_fd_sc_hd__xor2_1
  U1077
  (
    .A(A[9]),
    .B(n1233),
    .X(n1232)
  );


  sky130_fd_sc_hd__maj3_1
  U1078
  (
    .A(n1234),
    .B(n1235),
    .C(n1236),
    .X(n1230)
  );


  sky130_fd_sc_hd__xor2_1
  U1079
  (
    .A(A[9]),
    .B(n1237),
    .X(n1236)
  );


  sky130_fd_sc_hd__maj3_1
  U1080
  (
    .A(n1238),
    .B(n1239),
    .C(n1240),
    .X(n1234)
  );


  sky130_fd_sc_hd__xor2_1
  U1081
  (
    .A(A[9]),
    .B(n1241),
    .X(n1240)
  );


  sky130_fd_sc_hd__maj3_1
  U1082
  (
    .A(n1242),
    .B(n1243),
    .C(n1244),
    .X(n1238)
  );


  sky130_fd_sc_hd__xor2_1
  U1083
  (
    .A(A[9]),
    .B(n1245),
    .X(n1244)
  );


  sky130_fd_sc_hd__o22a_1
  U1084
  (
    .A1(n1246),
    .A2(n1247),
    .B1(n1246),
    .B2(n1248),
    .X(n1242)
  );


  sky130_fd_sc_hd__xnor2_1
  U1085
  (
    .A(n1249),
    .B(n408),
    .Y(n328)
  );


  sky130_fd_sc_hd__xnor2_1
  U1086
  (
    .A(n834),
    .B(n1174),
    .Y(n408)
  );


  sky130_fd_sc_hd__a221oi_1
  U1087
  (
    .A1(n1138),
    .A2(n807),
    .B1(n1139),
    .B2(n855),
    .C1(n1250),
    .Y(n1174)
  );


  sky130_fd_sc_hd__o22ai_1
  U1088
  (
    .A1(n815),
    .A2(n1022),
    .B1(n786),
    .B2(n1178),
    .Y(n1250)
  );


  sky130_fd_sc_hd__xnor2_1
  U1089
  (
    .A(n410),
    .B(n407),
    .Y(n1249)
  );


  sky130_fd_sc_hd__xnor2_1
  U1090
  (
    .A(n1145),
    .B(n1175),
    .Y(n407)
  );


  sky130_fd_sc_hd__a222oi_1
  U1091
  (
    .A1(n1251),
    .A2(n768),
    .B1(n1252),
    .B2(n741),
    .C1(n1253),
    .C2(n770),
    .Y(n1175)
  );


  sky130_fd_sc_hd__xnor2_1
  U1092
  (
    .A(n1254),
    .B(n1063),
    .Y(n410)
  );


  sky130_fd_sc_hd__xnor2_1
  U1093
  (
    .A(n1255),
    .B(n1196),
    .Y(n1063)
  );


  sky130_fd_sc_hd__xnor2_1
  U1094
  (
    .A(n751),
    .B(n1060),
    .Y(n1196)
  );


  sky130_fd_sc_hd__a221oi_1
  U1095
  (
    .A1(n861),
    .A2(B[9]),
    .B1(n1124),
    .B2(n862),
    .C1(n1256),
    .Y(n1060)
  );


  sky130_fd_sc_hd__o22ai_1
  U1096
  (
    .A1(n1029),
    .A2(n811),
    .B1(n970),
    .B2(n900),
    .Y(n1256)
  );


  sky130_fd_sc_hd__xnor2_1
  U1097
  (
    .A(n1195),
    .B(n1058),
    .Y(n1255)
  );


  sky130_fd_sc_hd__xnor2_1
  U1098
  (
    .A(n1257),
    .B(n951),
    .Y(n1058)
  );


  sky130_fd_sc_hd__xor2_1
  U1099
  (
    .A(n948),
    .B(n1258),
    .X(n951)
  );


  sky130_fd_sc_hd__xor2_1
  U1100
  (
    .A(A[15]),
    .B(n945),
    .X(n1258)
  );


  sky130_fd_sc_hd__clkinv_1
  U1101
  (
    .A(n949),
    .Y(n945)
  );


  sky130_fd_sc_hd__nand2_1
  U1102
  (
    .A(n740),
    .B(B[14]),
    .Y(n949)
  );


  sky130_fd_sc_hd__clkinv_1
  U1103
  (
    .A(n946),
    .Y(n948)
  );


  sky130_fd_sc_hd__xor2_1
  U1104
  (
    .A(n739),
    .B(n1259),
    .X(n946)
  );


  sky130_fd_sc_hd__a221oi_1
  U1105
  (
    .A1(n1260),
    .A2(n771),
    .B1(n767),
    .B2(B[13]),
    .C1(n1261),
    .Y(n1259)
  );


  sky130_fd_sc_hd__o22ai_1
  U1106
  (
    .A1(n1154),
    .A2(n809),
    .B1(n1262),
    .B2(n789),
    .Y(n1261)
  );


  sky130_fd_sc_hd__clkinv_1
  U1107
  (
    .A(n787),
    .Y(n767)
  );


  sky130_fd_sc_hd__xnor2_1
  U1108
  (
    .A(n1192),
    .B(n1191),
    .Y(n1257)
  );


  sky130_fd_sc_hd__o22ai_1
  U1109
  (
    .A1(n956),
    .A2(n957),
    .B1(n1263),
    .B2(n97),
    .Y(n1191)
  );


  sky130_fd_sc_hd__nor2_1
  U1110
  (
    .A(n953),
    .B(n954),
    .Y(n1263)
  );


  sky130_fd_sc_hd__o22ai_1
  U1111
  (
    .A1(n1264),
    .A2(n1265),
    .B1(n1266),
    .B2(n959),
    .Y(n1192)
  );


  sky130_fd_sc_hd__nor2_1
  U1112
  (
    .A(n1267),
    .B(n1268),
    .Y(n1266)
  );


  sky130_fd_sc_hd__clkinv_1
  U1113
  (
    .A(n1267),
    .Y(n1265)
  );


  sky130_fd_sc_hd__xnor2_1
  U1114
  (
    .A(n851),
    .B(n1061),
    .Y(n1195)
  );


  sky130_fd_sc_hd__a221oi_1
  U1115
  (
    .A1(n971),
    .A2(n982),
    .B1(n905),
    .B2(n980),
    .C1(n1269),
    .Y(n1061)
  );


  sky130_fd_sc_hd__o22ai_1
  U1116
  (
    .A1(n1003),
    .A2(n873),
    .B1(n1025),
    .B2(n876),
    .Y(n1269)
  );


  sky130_fd_sc_hd__xnor2_1
  U1117
  (
    .A(n1200),
    .B(n1199),
    .Y(n1254)
  );


  sky130_fd_sc_hd__o22ai_1
  U1118
  (
    .A1(n1270),
    .A2(n1271),
    .B1(n1272),
    .B2(n1066),
    .Y(n1199)
  );


  sky130_fd_sc_hd__and2_0
  U1119
  (
    .A(n1271),
    .B(n1270),
    .X(n1272)
  );


  sky130_fd_sc_hd__o22ai_1
  U1120
  (
    .A1(n1273),
    .A2(n1274),
    .B1(n1275),
    .B2(n1086),
    .Y(n1200)
  );


  sky130_fd_sc_hd__and2_0
  U1121
  (
    .A(n1274),
    .B(n1273),
    .X(n1275)
  );


  sky130_fd_sc_hd__maj3_1
  U1122
  (
    .A(n1276),
    .B(n318),
    .C(n1277),
    .X(n1201)
  );


  sky130_fd_sc_hd__maj3_1
  U1123
  (
    .A(n1278),
    .B(n418),
    .C(n1279),
    .X(n1277)
  );


  sky130_fd_sc_hd__xor2_1
  U1124
  (
    .A(A[12]),
    .B(n1280),
    .X(n1279)
  );


  sky130_fd_sc_hd__maj3_1
  U1125
  (
    .A(n1281),
    .B(n1282),
    .C(n1283),
    .X(n1278)
  );


  sky130_fd_sc_hd__xor2_1
  U1126
  (
    .A(A[12]),
    .B(n1284),
    .X(n1283)
  );


  sky130_fd_sc_hd__maj3_1
  U1127
  (
    .A(n1285),
    .B(n1286),
    .C(n1287),
    .X(n1281)
  );


  sky130_fd_sc_hd__xor2_1
  U1128
  (
    .A(A[12]),
    .B(n1288),
    .X(n1287)
  );


  sky130_fd_sc_hd__maj3_1
  U1129
  (
    .A(n1289),
    .B(n1290),
    .C(n1291),
    .X(n1285)
  );


  sky130_fd_sc_hd__xor2_1
  U1130
  (
    .A(A[12]),
    .B(n1292),
    .X(n1291)
  );


  sky130_fd_sc_hd__maj3_1
  U1131
  (
    .A(n1293),
    .B(n1294),
    .C(n1295),
    .X(n1289)
  );


  sky130_fd_sc_hd__xor2_1
  U1132
  (
    .A(A[12]),
    .B(n1296),
    .X(n1295)
  );


  sky130_fd_sc_hd__maj3_1
  U1133
  (
    .A(n1297),
    .B(n1298),
    .C(n1299),
    .X(n1293)
  );


  sky130_fd_sc_hd__xor2_1
  U1134
  (
    .A(A[12]),
    .B(n1300),
    .X(n1299)
  );


  sky130_fd_sc_hd__maj3_1
  U1135
  (
    .A(n1301),
    .B(n1302),
    .C(n1303),
    .X(n1297)
  );


  sky130_fd_sc_hd__xor2_1
  U1136
  (
    .A(A[12]),
    .B(n1304),
    .X(n1303)
  );


  sky130_fd_sc_hd__maj3_1
  U1137
  (
    .A(n1305),
    .B(n1306),
    .C(n1307),
    .X(n1301)
  );


  sky130_fd_sc_hd__xor2_1
  U1138
  (
    .A(A[12]),
    .B(n1308),
    .X(n1307)
  );


  sky130_fd_sc_hd__maj3_1
  U1139
  (
    .A(n1309),
    .B(n1310),
    .C(n1311),
    .X(n1305)
  );


  sky130_fd_sc_hd__xor2_1
  U1140
  (
    .A(A[12]),
    .B(n1312),
    .X(n1311)
  );


  sky130_fd_sc_hd__maj3_1
  U1141
  (
    .A(n1313),
    .B(n1314),
    .C(n1315),
    .X(n1309)
  );


  sky130_fd_sc_hd__xor2_1
  U1142
  (
    .A(A[12]),
    .B(n1316),
    .X(n1315)
  );


  sky130_fd_sc_hd__maj3_1
  U1143
  (
    .A(n1317),
    .B(n1318),
    .C(n1319),
    .X(n1313)
  );


  sky130_fd_sc_hd__xor2_1
  U1144
  (
    .A(A[12]),
    .B(n1320),
    .X(n1319)
  );


  sky130_fd_sc_hd__maj3_1
  U1145
  (
    .A(n1321),
    .B(n1322),
    .C(n1323),
    .X(n1317)
  );


  sky130_fd_sc_hd__xor2_1
  U1146
  (
    .A(A[12]),
    .B(n1324),
    .X(n1323)
  );


  sky130_fd_sc_hd__maj3_1
  U1147
  (
    .A(n1325),
    .B(n1326),
    .C(n1327),
    .X(n1321)
  );


  sky130_fd_sc_hd__xor2_1
  U1148
  (
    .A(A[12]),
    .B(n1328),
    .X(n1327)
  );


  sky130_fd_sc_hd__xnor2_1
  U1149
  (
    .A(n1329),
    .B(n454),
    .Y(n318)
  );


  sky130_fd_sc_hd__xnor2_1
  U1150
  (
    .A(n1330),
    .B(n1086),
    .Y(n454)
  );


  sky130_fd_sc_hd__xnor2_1
  U1151
  (
    .A(n1331),
    .B(n1066),
    .Y(n1086)
  );


  sky130_fd_sc_hd__xnor2_1
  U1152
  (
    .A(n1332),
    .B(n959),
    .Y(n1066)
  );


  sky130_fd_sc_hd__xor2_1
  U1153
  (
    .A(n956),
    .B(n1333),
    .X(n959)
  );


  sky130_fd_sc_hd__xor2_1
  U1154
  (
    .A(A[15]),
    .B(n953),
    .X(n1333)
  );


  sky130_fd_sc_hd__clkinv_1
  U1155
  (
    .A(n957),
    .Y(n953)
  );


  sky130_fd_sc_hd__nand2_1
  U1156
  (
    .A(n740),
    .B(B[15]),
    .Y(n957)
  );


  sky130_fd_sc_hd__clkinv_1
  U1157
  (
    .A(n954),
    .Y(n956)
  );


  sky130_fd_sc_hd__xor2_1
  U1158
  (
    .A(n739),
    .B(n1334),
    .X(n954)
  );


  sky130_fd_sc_hd__a221oi_1
  U1159
  (
    .A1(n769),
    .A2(B[13]),
    .B1(n783),
    .B2(B[12]),
    .C1(n1335),
    .Y(n1334)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1160
  (
    .B1(n1336),
    .B2(n787),
    .A1_N(n771),
    .A2_N(n1337),
    .Y(n1335)
  );


  sky130_fd_sc_hd__xor2_1
  U1161
  (
    .A(n1267),
    .B(n1264),
    .X(n1332)
  );


  sky130_fd_sc_hd__clkinv_1
  U1162
  (
    .A(n1268),
    .Y(n1264)
  );


  sky130_fd_sc_hd__o22ai_1
  U1163
  (
    .A1(n962),
    .A2(n1338),
    .B1(n1339),
    .B2(n963),
    .Y(n1268)
  );


  sky130_fd_sc_hd__and2_0
  U1164
  (
    .A(n1338),
    .B(n962),
    .X(n1339)
  );


  sky130_fd_sc_hd__xor2_1
  U1165
  (
    .A(n751),
    .B(n961),
    .X(n1267)
  );


  sky130_fd_sc_hd__a221oi_1
  U1166
  (
    .A1(n878),
    .A2(B[9]),
    .B1(n862),
    .B2(n1152),
    .C1(n1340),
    .Y(n961)
  );


  sky130_fd_sc_hd__o22ai_1
  U1167
  (
    .A1(n1154),
    .A2(n811),
    .B1(n1029),
    .B2(n880),
    .Y(n1340)
  );


  sky130_fd_sc_hd__xnor2_1
  U1168
  (
    .A(n1270),
    .B(n1271),
    .Y(n1331)
  );


  sky130_fd_sc_hd__xnor2_1
  U1169
  (
    .A(n851),
    .B(n1068),
    .Y(n1271)
  );


  sky130_fd_sc_hd__a221oi_1
  U1170
  (
    .A1(n905),
    .A2(n981),
    .B1(n995),
    .B2(n982),
    .C1(n1341),
    .Y(n1068)
  );


  sky130_fd_sc_hd__o22ai_1
  U1171
  (
    .A1(n901),
    .A2(n970),
    .B1(n1025),
    .B2(n873),
    .Y(n1341)
  );


  sky130_fd_sc_hd__o22a_1
  U1172
  (
    .A1(n1342),
    .A2(n1343),
    .B1(n1344),
    .B2(n1070),
    .X(n1270)
  );


  sky130_fd_sc_hd__and2_0
  U1173
  (
    .A(n1343),
    .B(n1342),
    .X(n1344)
  );


  sky130_fd_sc_hd__xnor2_1
  U1174
  (
    .A(n1273),
    .B(n1274),
    .Y(n1330)
  );


  sky130_fd_sc_hd__xnor2_1
  U1175
  (
    .A(n834),
    .B(n1088),
    .Y(n1274)
  );


  sky130_fd_sc_hd__a221oi_1
  U1176
  (
    .A1(n1164),
    .A2(n807),
    .B1(n1139),
    .B2(n874),
    .C1(n1345),
    .Y(n1088)
  );


  sky130_fd_sc_hd__o22ai_1
  U1177
  (
    .A1(n876),
    .A2(n1022),
    .B1(n815),
    .B2(n1166),
    .Y(n1345)
  );


  sky130_fd_sc_hd__o22a_1
  U1178
  (
    .A1(n1346),
    .A2(n1347),
    .B1(n1348),
    .B2(n1090),
    .X(n1273)
  );


  sky130_fd_sc_hd__and2_0
  U1179
  (
    .A(n1347),
    .B(n1346),
    .X(n1348)
  );


  sky130_fd_sc_hd__xnor2_1
  U1180
  (
    .A(n451),
    .B(n452),
    .Y(n1329)
  );


  sky130_fd_sc_hd__xnor2_1
  U1181
  (
    .A(n1145),
    .B(n1205),
    .Y(n452)
  );


  sky130_fd_sc_hd__a221oi_1
  U1182
  (
    .A1(n1349),
    .A2(n741),
    .B1(n1253),
    .B2(n784),
    .C1(n1350),
    .Y(n1205)
  );


  sky130_fd_sc_hd__o22ai_1
  U1183
  (
    .A1(n786),
    .A2(n1179),
    .B1(n788),
    .B2(n1351),
    .Y(n1350)
  );


  sky130_fd_sc_hd__o22a_1
  U1184
  (
    .A1(n1352),
    .A2(n1353),
    .B1(n1354),
    .B2(n1207),
    .X(n451)
  );


  sky130_fd_sc_hd__and2_0
  U1185
  (
    .A(n1353),
    .B(n1352),
    .X(n1354)
  );


  sky130_fd_sc_hd__maj3_1
  U1186
  (
    .A(n1355),
    .B(n311),
    .C(n1356),
    .X(n1276)
  );


  sky130_fd_sc_hd__xor2_1
  U1187
  (
    .A(n97),
    .B(n420),
    .X(n1356)
  );


  sky130_fd_sc_hd__o22ai_1
  U1188
  (
    .A1(n810),
    .A2(n1357),
    .B1(n813),
    .B2(n1358),
    .Y(n420)
  );


  sky130_fd_sc_hd__xnor2_1
  U1189
  (
    .A(n1359),
    .B(n418),
    .Y(n311)
  );


  sky130_fd_sc_hd__xnor2_1
  U1190
  (
    .A(n1360),
    .B(n1207),
    .Y(n418)
  );


  sky130_fd_sc_hd__xnor2_1
  U1191
  (
    .A(n1361),
    .B(n1090),
    .Y(n1207)
  );


  sky130_fd_sc_hd__xnor2_1
  U1192
  (
    .A(n1362),
    .B(n1070),
    .Y(n1090)
  );


  sky130_fd_sc_hd__xnor2_1
  U1193
  (
    .A(n1338),
    .B(n1363),
    .Y(n1070)
  );


  sky130_fd_sc_hd__xnor2_1
  U1194
  (
    .A(n963),
    .B(n962),
    .Y(n1363)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1195
  (
    .B1(n1364),
    .B2(n1365),
    .A1_N(n1366),
    .A2_N(n1367),
    .Y(n962)
  );


  sky130_fd_sc_hd__clkinv_1
  U1196
  (
    .A(n1365),
    .Y(n1366)
  );


  sky130_fd_sc_hd__nand2_1
  U1197
  (
    .A(n740),
    .B(B[16]),
    .Y(n963)
  );


  sky130_fd_sc_hd__xnor2_1
  U1198
  (
    .A(n739),
    .B(n965),
    .Y(n1338)
  );


  sky130_fd_sc_hd__a221oi_1
  U1199
  (
    .A1(n769),
    .A2(B[14]),
    .B1(n783),
    .B2(B[13]),
    .C1(n1368),
    .Y(n965)
  );


  sky130_fd_sc_hd__o22ai_1
  U1200
  (
    .A1(n1369),
    .A2(n787),
    .B1(n1370),
    .B2(n1371),
    .Y(n1368)
  );


  sky130_fd_sc_hd__xnor2_1
  U1201
  (
    .A(n1342),
    .B(n1343),
    .Y(n1362)
  );


  sky130_fd_sc_hd__xnor2_1
  U1202
  (
    .A(n751),
    .B(n1072),
    .Y(n1343)
  );


  sky130_fd_sc_hd__a221oi_1
  U1203
  (
    .A1(n862),
    .A2(n1187),
    .B1(n860),
    .B2(B[12]),
    .C1(n1372),
    .Y(n1072)
  );


  sky130_fd_sc_hd__o22ai_1
  U1204
  (
    .A1(n1029),
    .A2(n900),
    .B1(n1154),
    .B2(n880),
    .Y(n1372)
  );


  sky130_fd_sc_hd__o22a_1
  U1205
  (
    .A1(n1373),
    .A2(n1374),
    .B1(n1375),
    .B2(n1074),
    .X(n1342)
  );


  sky130_fd_sc_hd__and2_0
  U1206
  (
    .A(n1374),
    .B(n1373),
    .X(n1375)
  );


  sky130_fd_sc_hd__xnor2_1
  U1207
  (
    .A(n1346),
    .B(n1347),
    .Y(n1361)
  );


  sky130_fd_sc_hd__xnor2_1
  U1208
  (
    .A(n851),
    .B(n1092),
    .Y(n1347)
  );


  sky130_fd_sc_hd__a221oi_1
  U1209
  (
    .A1(n1035),
    .A2(n982),
    .B1(B[9]),
    .B2(n980),
    .C1(n1376),
    .Y(n1092)
  );


  sky130_fd_sc_hd__o22ai_1
  U1210
  (
    .A1(n1003),
    .A2(n970),
    .B1(n1025),
    .B2(n1037),
    .Y(n1376)
  );


  sky130_fd_sc_hd__o22a_1
  U1211
  (
    .A1(n1377),
    .A2(n1378),
    .B1(n1379),
    .B2(n1094),
    .X(n1346)
  );


  sky130_fd_sc_hd__and2_0
  U1212
  (
    .A(n1378),
    .B(n1377),
    .X(n1379)
  );


  sky130_fd_sc_hd__xnor2_1
  U1213
  (
    .A(n1352),
    .B(n1353),
    .Y(n1360)
  );


  sky130_fd_sc_hd__xnor2_1
  U1214
  (
    .A(n834),
    .B(n1209),
    .Y(n1353)
  );


  sky130_fd_sc_hd__a221oi_1
  U1215
  (
    .A1(n1139),
    .A2(n907),
    .B1(n1137),
    .B2(n908),
    .C1(n1380),
    .Y(n1209)
  );


  sky130_fd_sc_hd__o22ai_1
  U1216
  (
    .A1(n876),
    .A2(n1166),
    .B1(n815),
    .B2(n1178),
    .Y(n1380)
  );


  sky130_fd_sc_hd__o22a_1
  U1217
  (
    .A1(n1381),
    .A2(n1382),
    .B1(n1383),
    .B2(n1211),
    .X(n1352)
  );


  sky130_fd_sc_hd__and2_0
  U1218
  (
    .A(n1382),
    .B(n1381),
    .X(n1383)
  );


  sky130_fd_sc_hd__xnor2_1
  U1219
  (
    .A(n415),
    .B(n416),
    .Y(n1359)
  );


  sky130_fd_sc_hd__xnor2_1
  U1220
  (
    .A(n1145),
    .B(n1280),
    .Y(n416)
  );


  sky130_fd_sc_hd__a221oi_1
  U1221
  (
    .A1(n1253),
    .A2(n806),
    .B1(n1251),
    .B2(n807),
    .C1(n1384),
    .Y(n1280)
  );


  sky130_fd_sc_hd__o22ai_1
  U1222
  (
    .A1(n786),
    .A2(n1351),
    .B1(n788),
    .B2(n1385),
    .Y(n1384)
  );


  sky130_fd_sc_hd__o22a_1
  U1223
  (
    .A1(n1386),
    .A2(n1387),
    .B1(n1388),
    .B2(n1282),
    .X(n415)
  );


  sky130_fd_sc_hd__and2_0
  U1224
  (
    .A(n1387),
    .B(n1386),
    .X(n1388)
  );


  sky130_fd_sc_hd__maj3_1
  U1225
  (
    .A(n1389),
    .B(n304),
    .C(n1390),
    .X(n1355)
  );


  sky130_fd_sc_hd__xor2_1
  U1226
  (
    .A(A[15]),
    .B(n422),
    .X(n1390)
  );


  sky130_fd_sc_hd__a222oi_1
  U1227
  (
    .A1(n1391),
    .A2(n768),
    .B1(n1392),
    .B2(n741),
    .C1(n1393),
    .C2(n770),
    .Y(n422)
  );


  sky130_fd_sc_hd__xor2_1
  U1228
  (
    .A(n1394),
    .B(n741),
    .X(n770)
  );


  sky130_fd_sc_hd__xnor2_1
  U1229
  (
    .A(n1395),
    .B(n1282),
    .Y(n304)
  );


  sky130_fd_sc_hd__xnor2_1
  U1230
  (
    .A(n1396),
    .B(n1211),
    .Y(n1282)
  );


  sky130_fd_sc_hd__xnor2_1
  U1231
  (
    .A(n1397),
    .B(n1094),
    .Y(n1211)
  );


  sky130_fd_sc_hd__xnor2_1
  U1232
  (
    .A(n1398),
    .B(n1074),
    .Y(n1094)
  );


  sky130_fd_sc_hd__xor2_1
  U1233
  (
    .A(n1399),
    .B(n1365),
    .X(n1074)
  );


  sky130_fd_sc_hd__xor2_1
  U1234
  (
    .A(n739),
    .B(n1400),
    .X(n1365)
  );


  sky130_fd_sc_hd__a221oi_1
  U1235
  (
    .A1(n769),
    .A2(B[15]),
    .B1(n783),
    .B2(B[14]),
    .C1(n1401),
    .Y(n1400)
  );


  sky130_fd_sc_hd__o22ai_1
  U1236
  (
    .A1(n1402),
    .A2(n787),
    .B1(n1370),
    .B2(n1403),
    .Y(n1401)
  );


  sky130_fd_sc_hd__xor2_1
  U1237
  (
    .A(n1367),
    .B(n1364),
    .X(n1399)
  );


  sky130_fd_sc_hd__nor2_1
  U1238
  (
    .A(n1404),
    .B(n1405),
    .Y(n1364)
  );


  sky130_fd_sc_hd__nand2_1
  U1239
  (
    .A(n740),
    .B(B[17]),
    .Y(n1367)
  );


  sky130_fd_sc_hd__xnor2_1
  U1240
  (
    .A(n1373),
    .B(n1374),
    .Y(n1398)
  );


  sky130_fd_sc_hd__xnor2_1
  U1241
  (
    .A(n751),
    .B(n1076),
    .Y(n1374)
  );


  sky130_fd_sc_hd__a221oi_1
  U1242
  (
    .A1(n1260),
    .A2(n862),
    .B1(n860),
    .B2(B[13]),
    .C1(n1406),
    .Y(n1076)
  );


  sky130_fd_sc_hd__o22ai_1
  U1243
  (
    .A1(n1154),
    .A2(n900),
    .B1(n1262),
    .B2(n880),
    .Y(n1406)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1244
  (
    .B1(n1407),
    .B2(n1408),
    .A1_N(n1409),
    .A2_N(n1078),
    .Y(n1373)
  );


  sky130_fd_sc_hd__nor2_1
  U1245
  (
    .A(n1408),
    .B(n1407),
    .Y(n1409)
  );


  sky130_fd_sc_hd__xnor2_1
  U1246
  (
    .A(n1377),
    .B(n1378),
    .Y(n1397)
  );


  sky130_fd_sc_hd__xnor2_1
  U1247
  (
    .A(n851),
    .B(n1096),
    .Y(n1378)
  );


  sky130_fd_sc_hd__a221oi_1
  U1248
  (
    .A1(B[9]),
    .A2(n981),
    .B1(n1124),
    .B2(n982),
    .C1(n1410),
    .Y(n1096)
  );


  sky130_fd_sc_hd__o22ai_1
  U1249
  (
    .A1(n901),
    .A2(n1029),
    .B1(n1025),
    .B2(n970),
    .Y(n1410)
  );


  sky130_fd_sc_hd__o22a_1
  U1250
  (
    .A1(n1411),
    .A2(n1412),
    .B1(n1413),
    .B2(n1098),
    .X(n1377)
  );


  sky130_fd_sc_hd__and2_0
  U1251
  (
    .A(n1412),
    .B(n1411),
    .X(n1413)
  );


  sky130_fd_sc_hd__xnor2_1
  U1252
  (
    .A(n1381),
    .B(n1382),
    .Y(n1396)
  );


  sky130_fd_sc_hd__xnor2_1
  U1253
  (
    .A(n834),
    .B(n1213),
    .Y(n1382)
  );


  sky130_fd_sc_hd__a221oi_1
  U1254
  (
    .A1(n1139),
    .A2(n971),
    .B1(n1137),
    .B2(n905),
    .C1(n1414),
    .Y(n1213)
  );


  sky130_fd_sc_hd__o22ai_1
  U1255
  (
    .A1(n873),
    .A2(n1166),
    .B1(n876),
    .B2(n1178),
    .Y(n1414)
  );


  sky130_fd_sc_hd__o22a_1
  U1256
  (
    .A1(n1415),
    .A2(n1416),
    .B1(n1417),
    .B2(n1215),
    .X(n1381)
  );


  sky130_fd_sc_hd__and2_0
  U1257
  (
    .A(n1416),
    .B(n1415),
    .X(n1417)
  );


  sky130_fd_sc_hd__xnor2_1
  U1258
  (
    .A(n1386),
    .B(n1387),
    .Y(n1395)
  );


  sky130_fd_sc_hd__xnor2_1
  U1259
  (
    .A(n1145),
    .B(n1284),
    .Y(n1387)
  );


  sky130_fd_sc_hd__a221oi_1
  U1260
  (
    .A1(n1252),
    .A2(n807),
    .B1(n1253),
    .B2(n855),
    .C1(n1418),
    .Y(n1284)
  );


  sky130_fd_sc_hd__o22ai_1
  U1261
  (
    .A1(n815),
    .A2(n1179),
    .B1(n786),
    .B2(n1385),
    .Y(n1418)
  );


  sky130_fd_sc_hd__o22a_1
  U1262
  (
    .A1(n1419),
    .A2(n1420),
    .B1(n1421),
    .B2(n1286),
    .X(n1386)
  );


  sky130_fd_sc_hd__and2_0
  U1263
  (
    .A(n1420),
    .B(n1419),
    .X(n1421)
  );


  sky130_fd_sc_hd__maj3_1
  U1264
  (
    .A(n1422),
    .B(n297),
    .C(n1423),
    .X(n1389)
  );


  sky130_fd_sc_hd__xor2_1
  U1265
  (
    .A(A[15]),
    .B(n424),
    .X(n1423)
  );


  sky130_fd_sc_hd__a221oi_1
  U1266
  (
    .A1(n1424),
    .A2(n741),
    .B1(n1393),
    .B2(n784),
    .C1(n1425),
    .Y(n424)
  );


  sky130_fd_sc_hd__o22ai_1
  U1267
  (
    .A1(n786),
    .A2(n1357),
    .B1(n788),
    .B2(n1426),
    .Y(n1425)
  );


  sky130_fd_sc_hd__xnor2_1
  U1268
  (
    .A(n1427),
    .B(n1428),
    .Y(n784)
  );


  sky130_fd_sc_hd__xor2_1
  U1269
  (
    .A(n768),
    .B(n741),
    .X(n1428)
  );


  sky130_fd_sc_hd__xnor2_1
  U1270
  (
    .A(n1429),
    .B(n1286),
    .Y(n297)
  );


  sky130_fd_sc_hd__xnor2_1
  U1271
  (
    .A(n1430),
    .B(n1215),
    .Y(n1286)
  );


  sky130_fd_sc_hd__xnor2_1
  U1272
  (
    .A(n1431),
    .B(n1098),
    .Y(n1215)
  );


  sky130_fd_sc_hd__xnor2_1
  U1273
  (
    .A(n1432),
    .B(n1078),
    .Y(n1098)
  );


  sky130_fd_sc_hd__xnor2_1
  U1274
  (
    .A(n1404),
    .B(n1405),
    .Y(n1078)
  );


  sky130_fd_sc_hd__xnor2_1
  U1275
  (
    .A(n739),
    .B(n1433),
    .Y(n1405)
  );


  sky130_fd_sc_hd__a221oi_1
  U1276
  (
    .A1(n769),
    .A2(B[16]),
    .B1(n783),
    .B2(B[15]),
    .C1(n1434),
    .Y(n1433)
  );


  sky130_fd_sc_hd__o22ai_1
  U1277
  (
    .A1(n1435),
    .A2(n787),
    .B1(n1436),
    .B2(n1370),
    .Y(n1434)
  );


  sky130_fd_sc_hd__nand3_1
  U1278
  (
    .A(n740),
    .B(n1437),
    .C(n1438),
    .Y(n1404)
  );


  sky130_fd_sc_hd__xnor2_1
  U1279
  (
    .A(n1408),
    .B(n1407),
    .Y(n1432)
  );


  sky130_fd_sc_hd__o22ai_1
  U1280
  (
    .A1(n1081),
    .A2(n1439),
    .B1(n1440),
    .B2(n1082),
    .Y(n1407)
  );


  sky130_fd_sc_hd__and2_0
  U1281
  (
    .A(n1439),
    .B(n1081),
    .X(n1440)
  );


  sky130_fd_sc_hd__xnor2_1
  U1282
  (
    .A(n780),
    .B(n1080),
    .Y(n1408)
  );


  sky130_fd_sc_hd__a221oi_1
  U1283
  (
    .A1(n1337),
    .A2(n862),
    .B1(n860),
    .B2(B[14]),
    .C1(n1441),
    .Y(n1080)
  );


  sky130_fd_sc_hd__o22ai_1
  U1284
  (
    .A1(n1262),
    .A2(n900),
    .B1(n1185),
    .B2(n880),
    .Y(n1441)
  );


  sky130_fd_sc_hd__xnor2_1
  U1285
  (
    .A(n1411),
    .B(n1412),
    .Y(n1431)
  );


  sky130_fd_sc_hd__xnor2_1
  U1286
  (
    .A(n851),
    .B(n1100),
    .Y(n1412)
  );


  sky130_fd_sc_hd__a221oi_1
  U1287
  (
    .A1(B[9]),
    .A2(n1001),
    .B1(n1152),
    .B2(n982),
    .C1(n1442),
    .Y(n1100)
  );


  sky130_fd_sc_hd__o22ai_1
  U1288
  (
    .A1(n901),
    .A2(n1154),
    .B1(n1003),
    .B2(n1029),
    .Y(n1442)
  );


  sky130_fd_sc_hd__o22a_1
  U1289
  (
    .A1(n1443),
    .A2(n1444),
    .B1(n1445),
    .B2(n1102),
    .X(n1411)
  );


  sky130_fd_sc_hd__and2_0
  U1290
  (
    .A(n1444),
    .B(n1443),
    .X(n1445)
  );


  sky130_fd_sc_hd__xnor2_1
  U1291
  (
    .A(n1415),
    .B(n1416),
    .Y(n1430)
  );


  sky130_fd_sc_hd__xnor2_1
  U1292
  (
    .A(n834),
    .B(n1217),
    .Y(n1416)
  );


  sky130_fd_sc_hd__a221oi_1
  U1293
  (
    .A1(n1138),
    .A2(n905),
    .B1(n1139),
    .B2(n995),
    .C1(n1446),
    .Y(n1217)
  );


  sky130_fd_sc_hd__o22ai_1
  U1294
  (
    .A1(n970),
    .A2(n1022),
    .B1(n873),
    .B2(n1178),
    .Y(n1446)
  );


  sky130_fd_sc_hd__o22a_1
  U1295
  (
    .A1(n1447),
    .A2(n1448),
    .B1(n1449),
    .B2(n1219),
    .X(n1415)
  );


  sky130_fd_sc_hd__and2_0
  U1296
  (
    .A(n1448),
    .B(n1447),
    .X(n1449)
  );


  sky130_fd_sc_hd__xnor2_1
  U1297
  (
    .A(n1419),
    .B(n1420),
    .Y(n1429)
  );


  sky130_fd_sc_hd__xnor2_1
  U1298
  (
    .A(n1145),
    .B(n1288),
    .Y(n1420)
  );


  sky130_fd_sc_hd__a221oi_1
  U1299
  (
    .A1(n1349),
    .A2(n807),
    .B1(n1253),
    .B2(n874),
    .C1(n1450),
    .Y(n1288)
  );


  sky130_fd_sc_hd__o22ai_1
  U1300
  (
    .A1(n876),
    .A2(n1179),
    .B1(n815),
    .B2(n1351),
    .Y(n1450)
  );


  sky130_fd_sc_hd__o22a_1
  U1301
  (
    .A1(n1451),
    .A2(n1452),
    .B1(n1453),
    .B2(n1290),
    .X(n1419)
  );


  sky130_fd_sc_hd__and2_0
  U1302
  (
    .A(n1452),
    .B(n1451),
    .X(n1453)
  );


  sky130_fd_sc_hd__maj3_1
  U1303
  (
    .A(n1454),
    .B(n293),
    .C(n1455),
    .X(n1422)
  );


  sky130_fd_sc_hd__xor2_1
  U1304
  (
    .A(A[15]),
    .B(n426),
    .X(n1455)
  );


  sky130_fd_sc_hd__a221oi_1
  U1305
  (
    .A1(n1393),
    .A2(n806),
    .B1(n1391),
    .B2(n807),
    .C1(n1456),
    .Y(n426)
  );


  sky130_fd_sc_hd__o22ai_1
  U1306
  (
    .A1(n786),
    .A2(n1426),
    .B1(n788),
    .B2(n1457),
    .Y(n1456)
  );


  sky130_fd_sc_hd__xor2_1
  U1307
  (
    .A(n1458),
    .B(n1459),
    .X(n806)
  );


  sky130_fd_sc_hd__xor2_1
  U1308
  (
    .A(n768),
    .B(n1460),
    .X(n1459)
  );


  sky130_fd_sc_hd__xnor2_1
  U1309
  (
    .A(n1461),
    .B(n1290),
    .Y(n293)
  );


  sky130_fd_sc_hd__xnor2_1
  U1310
  (
    .A(n1462),
    .B(n1219),
    .Y(n1290)
  );


  sky130_fd_sc_hd__xnor2_1
  U1311
  (
    .A(n1463),
    .B(n1102),
    .Y(n1219)
  );


  sky130_fd_sc_hd__xnor2_1
  U1312
  (
    .A(n1464),
    .B(n1082),
    .Y(n1102)
  );


  sky130_fd_sc_hd__xnor2_1
  U1313
  (
    .A(n1438),
    .B(n1465),
    .Y(n1082)
  );


  sky130_fd_sc_hd__nor2b_1
  U1314
  (
    .B_N(n1437),
    .A(n739),
    .Y(n1465)
  );


  sky130_fd_sc_hd__xor2_1
  U1315
  (
    .A(n739),
    .B(n1466),
    .X(n1438)
  );


  sky130_fd_sc_hd__a222oi_1
  U1316
  (
    .A1(n771),
    .A2(n1467),
    .B1(n769),
    .B2(B[17]),
    .C1(n783),
    .C2(B[16]),
    .Y(n1466)
  );


  sky130_fd_sc_hd__clkinv_1
  U1317
  (
    .A(n789),
    .Y(n769)
  );


  sky130_fd_sc_hd__nand2_1
  U1318
  (
    .A(n1468),
    .B(n1469),
    .Y(n789)
  );


  sky130_fd_sc_hd__xnor2_1
  U1319
  (
    .A(n1439),
    .B(n1081),
    .Y(n1464)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1320
  (
    .B1(n1470),
    .B2(n1471),
    .A1_N(n1472),
    .A2_N(n1473),
    .Y(n1081)
  );


  sky130_fd_sc_hd__xnor2_1
  U1321
  (
    .A(n751),
    .B(n1084),
    .Y(n1439)
  );


  sky130_fd_sc_hd__a221oi_1
  U1322
  (
    .A1(n861),
    .A2(B[14]),
    .B1(n878),
    .B2(B[13]),
    .C1(n1474),
    .Y(n1084)
  );


  sky130_fd_sc_hd__o22ai_1
  U1323
  (
    .A1(n1369),
    .A2(n811),
    .B1(n812),
    .B2(n1371),
    .Y(n1474)
  );


  sky130_fd_sc_hd__xnor2_1
  U1324
  (
    .A(n1443),
    .B(n1444),
    .Y(n1463)
  );


  sky130_fd_sc_hd__xnor2_1
  U1325
  (
    .A(n851),
    .B(n1104),
    .Y(n1444)
  );


  sky130_fd_sc_hd__a221oi_1
  U1326
  (
    .A1(n1187),
    .A2(n982),
    .B1(B[12]),
    .B2(n980),
    .C1(n1475),
    .Y(n1104)
  );


  sky130_fd_sc_hd__o22ai_1
  U1327
  (
    .A1(n1025),
    .A2(n1029),
    .B1(n1003),
    .B2(n1154),
    .Y(n1475)
  );


  sky130_fd_sc_hd__o22a_1
  U1328
  (
    .A1(n1476),
    .A2(n1477),
    .B1(n1478),
    .B2(n1106),
    .X(n1443)
  );


  sky130_fd_sc_hd__and2_0
  U1329
  (
    .A(n1477),
    .B(n1476),
    .X(n1478)
  );


  sky130_fd_sc_hd__xnor2_1
  U1330
  (
    .A(n1447),
    .B(n1448),
    .Y(n1462)
  );


  sky130_fd_sc_hd__xnor2_1
  U1331
  (
    .A(n834),
    .B(n1221),
    .Y(n1448)
  );


  sky130_fd_sc_hd__a221oi_1
  U1332
  (
    .A1(n1139),
    .A2(n1035),
    .B1(n1137),
    .B2(B[9]),
    .C1(n1479),
    .Y(n1221)
  );


  sky130_fd_sc_hd__o22ai_1
  U1333
  (
    .A1(n970),
    .A2(n1166),
    .B1(n1037),
    .B2(n1178),
    .Y(n1479)
  );


  sky130_fd_sc_hd__o22a_1
  U1334
  (
    .A1(n1480),
    .A2(n1481),
    .B1(n1482),
    .B2(n1223),
    .X(n1447)
  );


  sky130_fd_sc_hd__and2_0
  U1335
  (
    .A(n1481),
    .B(n1480),
    .X(n1482)
  );


  sky130_fd_sc_hd__xnor2_1
  U1336
  (
    .A(n1451),
    .B(n1452),
    .Y(n1461)
  );


  sky130_fd_sc_hd__xnor2_1
  U1337
  (
    .A(n1145),
    .B(n1292),
    .Y(n1452)
  );


  sky130_fd_sc_hd__a221oi_1
  U1338
  (
    .A1(n1253),
    .A2(n907),
    .B1(n1251),
    .B2(n908),
    .C1(n1483),
    .Y(n1292)
  );


  sky130_fd_sc_hd__o22ai_1
  U1339
  (
    .A1(n876),
    .A2(n1351),
    .B1(n815),
    .B2(n1385),
    .Y(n1483)
  );


  sky130_fd_sc_hd__o22a_1
  U1340
  (
    .A1(n1484),
    .A2(n1485),
    .B1(n1486),
    .B2(n1294),
    .X(n1451)
  );


  sky130_fd_sc_hd__and2_0
  U1341
  (
    .A(n1485),
    .B(n1484),
    .X(n1486)
  );


  sky130_fd_sc_hd__maj3_1
  U1342
  (
    .A(n1487),
    .B(n159),
    .C(n1488),
    .X(n1454)
  );


  sky130_fd_sc_hd__xor2_1
  U1343
  (
    .A(A[15]),
    .B(n428),
    .X(n1488)
  );


  sky130_fd_sc_hd__a221oi_1
  U1344
  (
    .A1(n1392),
    .A2(n807),
    .B1(n1393),
    .B2(n855),
    .C1(n1489),
    .Y(n428)
  );


  sky130_fd_sc_hd__o22ai_1
  U1345
  (
    .A1(n815),
    .A2(n1357),
    .B1(n786),
    .B2(n1457),
    .Y(n1489)
  );


  sky130_fd_sc_hd__xor2_1
  U1346
  (
    .A(n1490),
    .B(n1491),
    .X(n855)
  );


  sky130_fd_sc_hd__xor2_1
  U1347
  (
    .A(n1460),
    .B(n807),
    .X(n1491)
  );


  sky130_fd_sc_hd__xnor2_1
  U1348
  (
    .A(n1492),
    .B(n1294),
    .Y(n159)
  );


  sky130_fd_sc_hd__xnor2_1
  U1349
  (
    .A(n1493),
    .B(n1223),
    .Y(n1294)
  );


  sky130_fd_sc_hd__xnor2_1
  U1350
  (
    .A(n1494),
    .B(n1106),
    .Y(n1223)
  );


  sky130_fd_sc_hd__xnor2_1
  U1351
  (
    .A(n1472),
    .B(n1495),
    .Y(n1106)
  );


  sky130_fd_sc_hd__xor2_1
  U1352
  (
    .A(n1470),
    .B(n1473),
    .X(n1495)
  );


  sky130_fd_sc_hd__clkinv_1
  U1353
  (
    .A(n1471),
    .Y(n1473)
  );


  sky130_fd_sc_hd__xor2_1
  U1354
  (
    .A(n751),
    .B(n1496),
    .X(n1471)
  );


  sky130_fd_sc_hd__a221oi_1
  U1355
  (
    .A1(n861),
    .A2(B[15]),
    .B1(n878),
    .B2(B[14]),
    .C1(n1497),
    .Y(n1496)
  );


  sky130_fd_sc_hd__o22ai_1
  U1356
  (
    .A1(n1402),
    .A2(n811),
    .B1(n812),
    .B2(n1403),
    .Y(n1497)
  );


  sky130_fd_sc_hd__nor2_1
  U1357
  (
    .A(n1498),
    .B(n1499),
    .Y(n1470)
  );


  sky130_fd_sc_hd__xor2_1
  U1358
  (
    .A(n1437),
    .B(n739),
    .X(n1472)
  );


  sky130_fd_sc_hd__xnor2_1
  U1359
  (
    .A(n739),
    .B(n1500),
    .Y(n1437)
  );


  sky130_fd_sc_hd__a21oi_1
  U1360
  (
    .A1(n1370),
    .A2(n809),
    .B1(n1435),
    .Y(n1500)
  );


  sky130_fd_sc_hd__clkinv_1
  U1361
  (
    .A(n783),
    .Y(n809)
  );


  sky130_fd_sc_hd__nor2_1
  U1362
  (
    .A(n1501),
    .B(n1468),
    .Y(n783)
  );


  sky130_fd_sc_hd__xnor2_1
  U1363
  (
    .A(n1476),
    .B(n1477),
    .Y(n1494)
  );


  sky130_fd_sc_hd__xnor2_1
  U1364
  (
    .A(n851),
    .B(n1108),
    .Y(n1477)
  );


  sky130_fd_sc_hd__a221oi_1
  U1365
  (
    .A1(n1260),
    .A2(n982),
    .B1(B[13]),
    .B2(n980),
    .C1(n1502),
    .Y(n1108)
  );


  sky130_fd_sc_hd__o22ai_1
  U1366
  (
    .A1(n1025),
    .A2(n1154),
    .B1(n1003),
    .B2(n1262),
    .Y(n1502)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1367
  (
    .B1(n1503),
    .B2(n1504),
    .A1_N(n1505),
    .A2_N(n1110),
    .Y(n1476)
  );


  sky130_fd_sc_hd__nor2_1
  U1368
  (
    .A(n1504),
    .B(n1503),
    .Y(n1505)
  );


  sky130_fd_sc_hd__xnor2_1
  U1369
  (
    .A(n1480),
    .B(n1481),
    .Y(n1493)
  );


  sky130_fd_sc_hd__xnor2_1
  U1370
  (
    .A(n834),
    .B(n1225),
    .Y(n1481)
  );


  sky130_fd_sc_hd__a221oi_1
  U1371
  (
    .A1(n1138),
    .A2(B[9]),
    .B1(n1139),
    .B2(n1124),
    .C1(n1506),
    .Y(n1225)
  );


  sky130_fd_sc_hd__o22ai_1
  U1372
  (
    .A1(n1029),
    .A2(n1022),
    .B1(n970),
    .B2(n1178),
    .Y(n1506)
  );


  sky130_fd_sc_hd__o22a_1
  U1373
  (
    .A1(n1507),
    .A2(n1508),
    .B1(n1509),
    .B2(n1227),
    .X(n1480)
  );


  sky130_fd_sc_hd__and2_0
  U1374
  (
    .A(n1508),
    .B(n1507),
    .X(n1509)
  );


  sky130_fd_sc_hd__xnor2_1
  U1375
  (
    .A(n1484),
    .B(n1485),
    .Y(n1492)
  );


  sky130_fd_sc_hd__xnor2_1
  U1376
  (
    .A(n1145),
    .B(n1296),
    .Y(n1485)
  );


  sky130_fd_sc_hd__a221oi_1
  U1377
  (
    .A1(n1253),
    .A2(n971),
    .B1(n1251),
    .B2(n905),
    .C1(n1510),
    .Y(n1296)
  );


  sky130_fd_sc_hd__o22ai_1
  U1378
  (
    .A1(n873),
    .A2(n1351),
    .B1(n876),
    .B2(n1385),
    .Y(n1510)
  );


  sky130_fd_sc_hd__o22a_1
  U1379
  (
    .A1(n1511),
    .A2(n1512),
    .B1(n1513),
    .B2(n1298),
    .X(n1484)
  );


  sky130_fd_sc_hd__and2_0
  U1380
  (
    .A(n1512),
    .B(n1511),
    .X(n1513)
  );


  sky130_fd_sc_hd__maj3_1
  U1381
  (
    .A(n1514),
    .B(n155),
    .C(n1515),
    .X(n1487)
  );


  sky130_fd_sc_hd__xor2_1
  U1382
  (
    .A(A[15]),
    .B(n430),
    .X(n1515)
  );


  sky130_fd_sc_hd__a221oi_1
  U1383
  (
    .A1(n1424),
    .A2(n807),
    .B1(n1393),
    .B2(n874),
    .C1(n1516),
    .Y(n430)
  );


  sky130_fd_sc_hd__o22ai_1
  U1384
  (
    .A1(n876),
    .A2(n1357),
    .B1(n815),
    .B2(n1426),
    .Y(n1516)
  );


  sky130_fd_sc_hd__xor2_1
  U1385
  (
    .A(n1517),
    .B(n1518),
    .X(n874)
  );


  sky130_fd_sc_hd__xor2_1
  U1386
  (
    .A(n807),
    .B(n1519),
    .X(n1518)
  );


  sky130_fd_sc_hd__xnor2_1
  U1387
  (
    .A(n1520),
    .B(n1298),
    .Y(n155)
  );


  sky130_fd_sc_hd__xnor2_1
  U1388
  (
    .A(n1521),
    .B(n1227),
    .Y(n1298)
  );


  sky130_fd_sc_hd__xnor2_1
  U1389
  (
    .A(n1522),
    .B(n1110),
    .Y(n1227)
  );


  sky130_fd_sc_hd__xnor2_1
  U1390
  (
    .A(n1498),
    .B(n1499),
    .Y(n1110)
  );


  sky130_fd_sc_hd__xnor2_1
  U1391
  (
    .A(n751),
    .B(n1523),
    .Y(n1499)
  );


  sky130_fd_sc_hd__a221oi_1
  U1392
  (
    .A1(n861),
    .A2(B[16]),
    .B1(n878),
    .B2(B[15]),
    .C1(n1524),
    .Y(n1523)
  );


  sky130_fd_sc_hd__o22ai_1
  U1393
  (
    .A1(n1435),
    .A2(n811),
    .B1(n1436),
    .B2(n812),
    .Y(n1524)
  );


  sky130_fd_sc_hd__clkinv_1
  U1394
  (
    .A(n860),
    .Y(n811)
  );


  sky130_fd_sc_hd__nor3b_1
  U1395
  (
    .C_N(n1525),
    .A(n1526),
    .B(n1527),
    .Y(n860)
  );


  sky130_fd_sc_hd__nand3_1
  U1396
  (
    .A(n780),
    .B(n1528),
    .C(n1529),
    .Y(n1498)
  );


  sky130_fd_sc_hd__clkinv_1
  U1397
  (
    .A(n751),
    .Y(n780)
  );


  sky130_fd_sc_hd__xnor2_1
  U1398
  (
    .A(n1504),
    .B(n1503),
    .Y(n1522)
  );


  sky130_fd_sc_hd__o22ai_1
  U1399
  (
    .A1(n1113),
    .A2(n1530),
    .B1(n1531),
    .B2(n1114),
    .Y(n1503)
  );


  sky130_fd_sc_hd__and2_0
  U1400
  (
    .A(n1530),
    .B(n1113),
    .X(n1531)
  );


  sky130_fd_sc_hd__xnor2_1
  U1401
  (
    .A(n872),
    .B(n1112),
    .Y(n1504)
  );


  sky130_fd_sc_hd__a221oi_1
  U1402
  (
    .A1(n1337),
    .A2(n982),
    .B1(B[14]),
    .B2(n980),
    .C1(n1532),
    .Y(n1112)
  );


  sky130_fd_sc_hd__o22ai_1
  U1403
  (
    .A1(n1025),
    .A2(n1262),
    .B1(n1003),
    .B2(n1185),
    .Y(n1532)
  );


  sky130_fd_sc_hd__clkinv_1
  U1404
  (
    .A(n901),
    .Y(n980)
  );


  sky130_fd_sc_hd__xnor2_1
  U1405
  (
    .A(n1507),
    .B(n1508),
    .Y(n1521)
  );


  sky130_fd_sc_hd__xnor2_1
  U1406
  (
    .A(n834),
    .B(n1229),
    .Y(n1508)
  );


  sky130_fd_sc_hd__a221oi_1
  U1407
  (
    .A1(n1164),
    .A2(B[9]),
    .B1(n1139),
    .B2(n1152),
    .C1(n1533),
    .Y(n1229)
  );


  sky130_fd_sc_hd__o22ai_1
  U1408
  (
    .A1(n1154),
    .A2(n1022),
    .B1(n1029),
    .B2(n1166),
    .Y(n1533)
  );


  sky130_fd_sc_hd__o22a_1
  U1409
  (
    .A1(n1534),
    .A2(n1535),
    .B1(n1536),
    .B2(n1231),
    .X(n1507)
  );


  sky130_fd_sc_hd__and2_0
  U1410
  (
    .A(n1535),
    .B(n1534),
    .X(n1536)
  );


  sky130_fd_sc_hd__xnor2_1
  U1411
  (
    .A(n1511),
    .B(n1512),
    .Y(n1520)
  );


  sky130_fd_sc_hd__xnor2_1
  U1412
  (
    .A(n1145),
    .B(n1300),
    .Y(n1512)
  );


  sky130_fd_sc_hd__a221oi_1
  U1413
  (
    .A1(n1252),
    .A2(n905),
    .B1(n1253),
    .B2(n995),
    .C1(n1537),
    .Y(n1300)
  );


  sky130_fd_sc_hd__o22ai_1
  U1414
  (
    .A1(n970),
    .A2(n1179),
    .B1(n873),
    .B2(n1385),
    .Y(n1537)
  );


  sky130_fd_sc_hd__o22a_1
  U1415
  (
    .A1(n1538),
    .A2(n1539),
    .B1(n1540),
    .B2(n1302),
    .X(n1511)
  );


  sky130_fd_sc_hd__and2_0
  U1416
  (
    .A(n1539),
    .B(n1538),
    .X(n1540)
  );


  sky130_fd_sc_hd__maj3_1
  U1417
  (
    .A(n1541),
    .B(n151),
    .C(n1542),
    .X(n1514)
  );


  sky130_fd_sc_hd__xor2_1
  U1418
  (
    .A(A[15]),
    .B(n432),
    .X(n1542)
  );


  sky130_fd_sc_hd__a221oi_1
  U1419
  (
    .A1(n1393),
    .A2(n907),
    .B1(n1391),
    .B2(n908),
    .C1(n1543),
    .Y(n432)
  );


  sky130_fd_sc_hd__o22ai_1
  U1420
  (
    .A1(n876),
    .A2(n1426),
    .B1(n815),
    .B2(n1457),
    .Y(n1543)
  );


  sky130_fd_sc_hd__xor2_1
  U1421
  (
    .A(n1544),
    .B(n1545),
    .X(n907)
  );


  sky130_fd_sc_hd__xor2_1
  U1422
  (
    .A(n1519),
    .B(n853),
    .X(n1545)
  );


  sky130_fd_sc_hd__xnor2_1
  U1423
  (
    .A(n1546),
    .B(n1302),
    .Y(n151)
  );


  sky130_fd_sc_hd__xnor2_1
  U1424
  (
    .A(n1547),
    .B(n1231),
    .Y(n1302)
  );


  sky130_fd_sc_hd__xnor2_1
  U1425
  (
    .A(n1548),
    .B(n1114),
    .Y(n1231)
  );


  sky130_fd_sc_hd__xnor2_1
  U1426
  (
    .A(n1529),
    .B(n1549),
    .Y(n1114)
  );


  sky130_fd_sc_hd__nor2b_1
  U1427
  (
    .B_N(n1528),
    .A(n751),
    .Y(n1549)
  );


  sky130_fd_sc_hd__xor2_1
  U1428
  (
    .A(n751),
    .B(n1550),
    .X(n1529)
  );


  sky130_fd_sc_hd__a222oi_1
  U1429
  (
    .A1(n862),
    .A2(n1467),
    .B1(n861),
    .B2(B[17]),
    .C1(n878),
    .C2(B[16]),
    .Y(n1550)
  );


  sky130_fd_sc_hd__clkinv_1
  U1430
  (
    .A(n880),
    .Y(n861)
  );


  sky130_fd_sc_hd__nand2_1
  U1431
  (
    .A(n1551),
    .B(n1526),
    .Y(n880)
  );


  sky130_fd_sc_hd__xor2_1
  U1432
  (
    .A(n1552),
    .B(n1553),
    .X(n1526)
  );


  sky130_fd_sc_hd__clkinv_1
  U1433
  (
    .A(n812),
    .Y(n862)
  );


  sky130_fd_sc_hd__xnor2_1
  U1434
  (
    .A(n1530),
    .B(n1113),
    .Y(n1548)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1435
  (
    .B1(n1554),
    .B2(n1555),
    .A1_N(n1556),
    .A2_N(n1557),
    .Y(n1113)
  );


  sky130_fd_sc_hd__xnor2_1
  U1436
  (
    .A(n851),
    .B(n1116),
    .Y(n1530)
  );


  sky130_fd_sc_hd__a221oi_1
  U1437
  (
    .A1(B[14]),
    .A2(n981),
    .B1(B[13]),
    .B2(n1001),
    .C1(n1558),
    .Y(n1116)
  );


  sky130_fd_sc_hd__o22ai_1
  U1438
  (
    .A1(n901),
    .A2(n1369),
    .B1(n902),
    .B2(n1371),
    .Y(n1558)
  );


  sky130_fd_sc_hd__clkinv_1
  U1439
  (
    .A(n1559),
    .Y(n1371)
  );


  sky130_fd_sc_hd__xnor2_1
  U1440
  (
    .A(n1534),
    .B(n1535),
    .Y(n1547)
  );


  sky130_fd_sc_hd__xnor2_1
  U1441
  (
    .A(n834),
    .B(n1233),
    .Y(n1535)
  );


  sky130_fd_sc_hd__a221oi_1
  U1442
  (
    .A1(n1139),
    .A2(n1187),
    .B1(n1137),
    .B2(B[12]),
    .C1(n1560),
    .Y(n1233)
  );


  sky130_fd_sc_hd__o22ai_1
  U1443
  (
    .A1(n1029),
    .A2(n1178),
    .B1(n1154),
    .B2(n1166),
    .Y(n1560)
  );


  sky130_fd_sc_hd__o22a_1
  U1444
  (
    .A1(n1561),
    .A2(n1562),
    .B1(n1563),
    .B2(n1235),
    .X(n1534)
  );


  sky130_fd_sc_hd__and2_0
  U1445
  (
    .A(n1562),
    .B(n1561),
    .X(n1563)
  );


  sky130_fd_sc_hd__xnor2_1
  U1446
  (
    .A(n1538),
    .B(n1539),
    .Y(n1546)
  );


  sky130_fd_sc_hd__xnor2_1
  U1447
  (
    .A(n1145),
    .B(n1304),
    .Y(n1539)
  );


  sky130_fd_sc_hd__a221oi_1
  U1448
  (
    .A1(n1253),
    .A2(n1035),
    .B1(n1251),
    .B2(B[9]),
    .C1(n1564),
    .Y(n1304)
  );


  sky130_fd_sc_hd__o22ai_1
  U1449
  (
    .A1(n970),
    .A2(n1351),
    .B1(n1037),
    .B2(n1385),
    .Y(n1564)
  );


  sky130_fd_sc_hd__o22a_1
  U1450
  (
    .A1(n1565),
    .A2(n1566),
    .B1(n1567),
    .B2(n1306),
    .X(n1538)
  );


  sky130_fd_sc_hd__and2_0
  U1451
  (
    .A(n1566),
    .B(n1565),
    .X(n1567)
  );


  sky130_fd_sc_hd__maj3_1
  U1452
  (
    .A(n1568),
    .B(n147),
    .C(n1569),
    .X(n1541)
  );


  sky130_fd_sc_hd__xor2_1
  U1453
  (
    .A(A[15]),
    .B(n434),
    .X(n1569)
  );


  sky130_fd_sc_hd__a221oi_1
  U1454
  (
    .A1(n1393),
    .A2(n971),
    .B1(n1391),
    .B2(n905),
    .C1(n1570),
    .Y(n434)
  );


  sky130_fd_sc_hd__o22ai_1
  U1455
  (
    .A1(n873),
    .A2(n1426),
    .B1(n876),
    .B2(n1457),
    .Y(n1570)
  );


  sky130_fd_sc_hd__xnor2_1
  U1456
  (
    .A(n1571),
    .B(n1572),
    .Y(n971)
  );


  sky130_fd_sc_hd__xor2_1
  U1457
  (
    .A(n853),
    .B(n908),
    .X(n1572)
  );


  sky130_fd_sc_hd__xnor2_1
  U1458
  (
    .A(n1573),
    .B(n1306),
    .Y(n147)
  );


  sky130_fd_sc_hd__xnor2_1
  U1459
  (
    .A(n1574),
    .B(n1235),
    .Y(n1306)
  );


  sky130_fd_sc_hd__xnor2_1
  U1460
  (
    .A(n1556),
    .B(n1575),
    .Y(n1235)
  );


  sky130_fd_sc_hd__xor2_1
  U1461
  (
    .A(n1554),
    .B(n1557),
    .X(n1575)
  );


  sky130_fd_sc_hd__clkinv_1
  U1462
  (
    .A(n1555),
    .Y(n1557)
  );


  sky130_fd_sc_hd__xor2_1
  U1463
  (
    .A(n851),
    .B(n1576),
    .X(n1555)
  );


  sky130_fd_sc_hd__a221oi_1
  U1464
  (
    .A1(B[15]),
    .A2(n981),
    .B1(B[14]),
    .B2(n1001),
    .C1(n1577),
    .Y(n1576)
  );


  sky130_fd_sc_hd__o22ai_1
  U1465
  (
    .A1(n901),
    .A2(n1402),
    .B1(n902),
    .B2(n1403),
    .Y(n1577)
  );


  sky130_fd_sc_hd__nor2_1
  U1466
  (
    .A(n1578),
    .B(n1579),
    .Y(n1554)
  );


  sky130_fd_sc_hd__xor2_1
  U1467
  (
    .A(n1528),
    .B(n751),
    .X(n1556)
  );


  sky130_fd_sc_hd__xnor2_1
  U1468
  (
    .A(n751),
    .B(n1580),
    .Y(n1528)
  );


  sky130_fd_sc_hd__a21oi_1
  U1469
  (
    .A1(n812),
    .A2(n900),
    .B1(n1435),
    .Y(n1580)
  );


  sky130_fd_sc_hd__clkinv_1
  U1470
  (
    .A(n878),
    .Y(n900)
  );


  sky130_fd_sc_hd__nor2_1
  U1471
  (
    .A(n1525),
    .B(n1551),
    .Y(n878)
  );


  sky130_fd_sc_hd__clkinv_1
  U1472
  (
    .A(n1527),
    .Y(n1551)
  );


  sky130_fd_sc_hd__nand2_1
  U1473
  (
    .A(n1527),
    .B(n1525),
    .Y(n812)
  );


  sky130_fd_sc_hd__xnor2_1
  U1474
  (
    .A(n751),
    .B(n1552),
    .Y(n1525)
  );


  sky130_fd_sc_hd__nor2_1
  U1475
  (
    .A(n720),
    .B(MODE_0_0),
    .Y(n1552)
  );


  sky130_fd_sc_hd__clkinv_1
  U1476
  (
    .A(A[4]),
    .Y(n720)
  );


  sky130_fd_sc_hd__xor2_1
  U1477
  (
    .A(n1553),
    .B(n872),
    .X(n1527)
  );


  sky130_fd_sc_hd__nor2_1
  U1478
  (
    .A(n515),
    .B(MODE_0_0),
    .Y(n1553)
  );


  sky130_fd_sc_hd__clkinv_1
  U1479
  (
    .A(A[5]),
    .Y(n515)
  );


  sky130_fd_sc_hd__xnor2_1
  U1480
  (
    .A(n1561),
    .B(n1562),
    .Y(n1574)
  );


  sky130_fd_sc_hd__xnor2_1
  U1481
  (
    .A(n834),
    .B(n1237),
    .Y(n1562)
  );


  sky130_fd_sc_hd__a221oi_1
  U1482
  (
    .A1(n1139),
    .A2(n1260),
    .B1(n1137),
    .B2(B[13]),
    .C1(n1581),
    .Y(n1237)
  );


  sky130_fd_sc_hd__o22ai_1
  U1483
  (
    .A1(n1154),
    .A2(n1178),
    .B1(n1262),
    .B2(n1166),
    .Y(n1581)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1484
  (
    .B1(n1582),
    .B2(n1583),
    .A1_N(n1584),
    .A2_N(n1239),
    .Y(n1561)
  );


  sky130_fd_sc_hd__nor2_1
  U1485
  (
    .A(n1583),
    .B(n1582),
    .Y(n1584)
  );


  sky130_fd_sc_hd__xnor2_1
  U1486
  (
    .A(n1565),
    .B(n1566),
    .Y(n1573)
  );


  sky130_fd_sc_hd__xnor2_1
  U1487
  (
    .A(n1145),
    .B(n1308),
    .Y(n1566)
  );


  sky130_fd_sc_hd__a221oi_1
  U1488
  (
    .A1(n1252),
    .A2(B[9]),
    .B1(n1253),
    .B2(n1124),
    .C1(n1585),
    .Y(n1308)
  );


  sky130_fd_sc_hd__o22ai_1
  U1489
  (
    .A1(n1029),
    .A2(n1179),
    .B1(n970),
    .B2(n1385),
    .Y(n1585)
  );


  sky130_fd_sc_hd__o22a_1
  U1490
  (
    .A1(n1586),
    .A2(n1587),
    .B1(n1588),
    .B2(n1310),
    .X(n1565)
  );


  sky130_fd_sc_hd__and2_0
  U1491
  (
    .A(n1587),
    .B(n1586),
    .X(n1588)
  );


  sky130_fd_sc_hd__maj3_1
  U1492
  (
    .A(n1589),
    .B(n143),
    .C(n1590),
    .X(n1568)
  );


  sky130_fd_sc_hd__xor2_1
  U1493
  (
    .A(A[15]),
    .B(n436),
    .X(n1590)
  );


  sky130_fd_sc_hd__a221oi_1
  U1494
  (
    .A1(n1392),
    .A2(n905),
    .B1(n1393),
    .B2(n995),
    .C1(n1591),
    .Y(n436)
  );


  sky130_fd_sc_hd__o22ai_1
  U1495
  (
    .A1(n970),
    .A2(n1357),
    .B1(n873),
    .B2(n1457),
    .Y(n1591)
  );


  sky130_fd_sc_hd__xor2_1
  U1496
  (
    .A(n1592),
    .B(n1593),
    .X(n995)
  );


  sky130_fd_sc_hd__xor2_1
  U1497
  (
    .A(n908),
    .B(n905),
    .X(n1593)
  );


  sky130_fd_sc_hd__xnor2_1
  U1498
  (
    .A(n1594),
    .B(n1310),
    .Y(n143)
  );


  sky130_fd_sc_hd__xor2_1
  U1499
  (
    .A(n1239),
    .B(n1595),
    .X(n1310)
  );


  sky130_fd_sc_hd__xor2_1
  U1500
  (
    .A(n1582),
    .B(n1583),
    .X(n1595)
  );


  sky130_fd_sc_hd__xor2_1
  U1501
  (
    .A(n834),
    .B(n1241),
    .X(n1583)
  );


  sky130_fd_sc_hd__a221oi_1
  U1502
  (
    .A1(n1139),
    .A2(n1337),
    .B1(n1137),
    .B2(B[14]),
    .C1(n1596),
    .Y(n1241)
  );


  sky130_fd_sc_hd__o22ai_1
  U1503
  (
    .A1(n1262),
    .A2(n1178),
    .B1(n1185),
    .B2(n1166),
    .Y(n1596)
  );


  sky130_fd_sc_hd__o22ai_1
  U1504
  (
    .A1(n1597),
    .A2(n1598),
    .B1(n1599),
    .B2(n1243),
    .Y(n1582)
  );


  sky130_fd_sc_hd__nor2_1
  U1505
  (
    .A(n1600),
    .B(n1601),
    .Y(n1599)
  );


  sky130_fd_sc_hd__clkinv_1
  U1506
  (
    .A(n1600),
    .Y(n1598)
  );


  sky130_fd_sc_hd__xnor2_1
  U1507
  (
    .A(n1578),
    .B(n1579),
    .Y(n1239)
  );


  sky130_fd_sc_hd__xnor2_1
  U1508
  (
    .A(n851),
    .B(n1602),
    .Y(n1579)
  );


  sky130_fd_sc_hd__a221oi_1
  U1509
  (
    .A1(B[16]),
    .A2(n981),
    .B1(B[15]),
    .B2(n1001),
    .C1(n1603),
    .Y(n1602)
  );


  sky130_fd_sc_hd__o22ai_1
  U1510
  (
    .A1(n901),
    .A2(n1435),
    .B1(n1436),
    .B2(n902),
    .Y(n1603)
  );


  sky130_fd_sc_hd__nand3_1
  U1511
  (
    .A(n1604),
    .B(n1605),
    .C(n1606),
    .Y(n901)
  );


  sky130_fd_sc_hd__nand3_1
  U1512
  (
    .A(n872),
    .B(n1607),
    .C(n1608),
    .Y(n1578)
  );


  sky130_fd_sc_hd__xnor2_1
  U1513
  (
    .A(n1586),
    .B(n1587),
    .Y(n1594)
  );


  sky130_fd_sc_hd__xnor2_1
  U1514
  (
    .A(n1145),
    .B(n1312),
    .Y(n1587)
  );


  sky130_fd_sc_hd__a221oi_1
  U1515
  (
    .A1(n1349),
    .A2(B[9]),
    .B1(n1253),
    .B2(n1152),
    .C1(n1609),
    .Y(n1312)
  );


  sky130_fd_sc_hd__o22ai_1
  U1516
  (
    .A1(n1154),
    .A2(n1179),
    .B1(n1029),
    .B2(n1351),
    .Y(n1609)
  );


  sky130_fd_sc_hd__o22a_1
  U1517
  (
    .A1(n1610),
    .A2(n1611),
    .B1(n1612),
    .B2(n1314),
    .X(n1586)
  );


  sky130_fd_sc_hd__and2_0
  U1518
  (
    .A(n1611),
    .B(n1610),
    .X(n1612)
  );


  sky130_fd_sc_hd__maj3_1
  U1519
  (
    .A(n1613),
    .B(n139),
    .C(n1614),
    .X(n1589)
  );


  sky130_fd_sc_hd__xor2_1
  U1520
  (
    .A(A[15]),
    .B(n438),
    .X(n1614)
  );


  sky130_fd_sc_hd__a221oi_1
  U1521
  (
    .A1(n1393),
    .A2(n1035),
    .B1(n1391),
    .B2(B[9]),
    .C1(n1615),
    .Y(n438)
  );


  sky130_fd_sc_hd__o22ai_1
  U1522
  (
    .A1(n970),
    .A2(n1426),
    .B1(n1037),
    .B2(n1457),
    .Y(n1615)
  );


  sky130_fd_sc_hd__xor2_1
  U1523
  (
    .A(n1616),
    .B(n1617),
    .X(n1035)
  );


  sky130_fd_sc_hd__xor2_1
  U1524
  (
    .A(n1037),
    .B(n970),
    .X(n1617)
  );


  sky130_fd_sc_hd__xnor2_1
  U1525
  (
    .A(n1618),
    .B(n1314),
    .Y(n139)
  );


  sky130_fd_sc_hd__xnor2_1
  U1526
  (
    .A(n1619),
    .B(n1243),
    .Y(n1314)
  );


  sky130_fd_sc_hd__xnor2_1
  U1527
  (
    .A(n1608),
    .B(n1620),
    .Y(n1243)
  );


  sky130_fd_sc_hd__nor2b_1
  U1528
  (
    .B_N(n1607),
    .A(n851),
    .Y(n1620)
  );


  sky130_fd_sc_hd__xor2_1
  U1529
  (
    .A(n851),
    .B(n1621),
    .X(n1608)
  );


  sky130_fd_sc_hd__a222oi_1
  U1530
  (
    .A1(n982),
    .A2(n1467),
    .B1(B[17]),
    .B2(n981),
    .C1(B[16]),
    .C2(n1001),
    .Y(n1621)
  );


  sky130_fd_sc_hd__clkinv_1
  U1531
  (
    .A(n1025),
    .Y(n1001)
  );


  sky130_fd_sc_hd__clkinv_1
  U1532
  (
    .A(n1003),
    .Y(n981)
  );


  sky130_fd_sc_hd__nand2_1
  U1533
  (
    .A(n1604),
    .B(n1622),
    .Y(n1003)
  );


  sky130_fd_sc_hd__clkinv_1
  U1534
  (
    .A(n1606),
    .Y(n1622)
  );


  sky130_fd_sc_hd__xor2_1
  U1535
  (
    .A(n1623),
    .B(n1624),
    .X(n1606)
  );


  sky130_fd_sc_hd__clkinv_1
  U1536
  (
    .A(n902),
    .Y(n982)
  );


  sky130_fd_sc_hd__xor2_1
  U1537
  (
    .A(n1600),
    .B(n1597),
    .X(n1619)
  );


  sky130_fd_sc_hd__clkinv_1
  U1538
  (
    .A(n1601),
    .Y(n1597)
  );


  sky130_fd_sc_hd__o22ai_1
  U1539
  (
    .A1(n1246),
    .A2(n1248),
    .B1(n1247),
    .B2(n1246),
    .Y(n1601)
  );


  sky130_fd_sc_hd__xor2_1
  U1540
  (
    .A(n834),
    .B(n1245),
    .X(n1600)
  );


  sky130_fd_sc_hd__a221oi_1
  U1541
  (
    .A1(n1139),
    .A2(n1559),
    .B1(n1137),
    .B2(B[15]),
    .C1(n1625),
    .Y(n1245)
  );


  sky130_fd_sc_hd__o22ai_1
  U1542
  (
    .A1(n1185),
    .A2(n1178),
    .B1(n1336),
    .B2(n1166),
    .Y(n1625)
  );


  sky130_fd_sc_hd__xnor2_1
  U1543
  (
    .A(n1610),
    .B(n1611),
    .Y(n1618)
  );


  sky130_fd_sc_hd__xnor2_1
  U1544
  (
    .A(n1145),
    .B(n1316),
    .Y(n1611)
  );


  sky130_fd_sc_hd__a221oi_1
  U1545
  (
    .A1(n1253),
    .A2(n1187),
    .B1(n1251),
    .B2(B[12]),
    .C1(n1626),
    .Y(n1316)
  );


  sky130_fd_sc_hd__o22ai_1
  U1546
  (
    .A1(n1029),
    .A2(n1385),
    .B1(n1154),
    .B2(n1351),
    .Y(n1626)
  );


  sky130_fd_sc_hd__o22a_1
  U1547
  (
    .A1(n1627),
    .A2(n1628),
    .B1(n1629),
    .B2(n1318),
    .X(n1610)
  );


  sky130_fd_sc_hd__and2_0
  U1548
  (
    .A(n1628),
    .B(n1627),
    .X(n1629)
  );


  sky130_fd_sc_hd__maj3_1
  U1549
  (
    .A(n1630),
    .B(n135),
    .C(n1631),
    .X(n1613)
  );


  sky130_fd_sc_hd__xor2_1
  U1550
  (
    .A(A[15]),
    .B(n440),
    .X(n1631)
  );


  sky130_fd_sc_hd__a221oi_1
  U1551
  (
    .A1(n1392),
    .A2(B[9]),
    .B1(n1393),
    .B2(n1124),
    .C1(n1632),
    .Y(n440)
  );


  sky130_fd_sc_hd__o22ai_1
  U1552
  (
    .A1(n1029),
    .A2(n1357),
    .B1(n970),
    .B2(n1457),
    .Y(n1632)
  );


  sky130_fd_sc_hd__xor2_1
  U1553
  (
    .A(n1633),
    .B(n1634),
    .X(n1124)
  );


  sky130_fd_sc_hd__xor2_1
  U1554
  (
    .A(n993),
    .B(n970),
    .X(n1634)
  );


  sky130_fd_sc_hd__xnor2_1
  U1555
  (
    .A(n1635),
    .B(n1318),
    .Y(n135)
  );


  sky130_fd_sc_hd__xnor2_1
  U1556
  (
    .A(n1247),
    .B(n1636),
    .Y(n1318)
  );


  sky130_fd_sc_hd__xnor2_1
  U1557
  (
    .A(n1248),
    .B(n1246),
    .Y(n1636)
  );


  sky130_fd_sc_hd__xnor2_1
  U1558
  (
    .A(n834),
    .B(n1637),
    .Y(n1246)
  );


  sky130_fd_sc_hd__a221oi_1
  U1559
  (
    .A1(n1139),
    .A2(n1638),
    .B1(n1137),
    .B2(B[16]),
    .C1(n1639),
    .Y(n1637)
  );


  sky130_fd_sc_hd__o22ai_1
  U1560
  (
    .A1(n1336),
    .A2(n1178),
    .B1(n1369),
    .B2(n1166),
    .Y(n1639)
  );


  sky130_fd_sc_hd__or2_0
  U1561
  (
    .A(n1640),
    .B(n1641),
    .X(n1248)
  );


  sky130_fd_sc_hd__xor2_1
  U1562
  (
    .A(n1607),
    .B(n851),
    .X(n1247)
  );


  sky130_fd_sc_hd__xnor2_1
  U1563
  (
    .A(n851),
    .B(n1642),
    .Y(n1607)
  );


  sky130_fd_sc_hd__a21oi_1
  U1564
  (
    .A1(n902),
    .A2(n1025),
    .B1(n1435),
    .Y(n1642)
  );


  sky130_fd_sc_hd__nand2_1
  U1565
  (
    .A(n1643),
    .B(n1644),
    .Y(n1025)
  );


  sky130_fd_sc_hd__nand2_1
  U1566
  (
    .A(n1605),
    .B(n1644),
    .Y(n902)
  );


  sky130_fd_sc_hd__clkinv_1
  U1567
  (
    .A(n1604),
    .Y(n1644)
  );


  sky130_fd_sc_hd__xor2_1
  U1568
  (
    .A(n834),
    .B(n1624),
    .X(n1604)
  );


  sky130_fd_sc_hd__nor2_1
  U1569
  (
    .A(n301),
    .B(MODE_0_0),
    .Y(n1624)
  );


  sky130_fd_sc_hd__clkinv_1
  U1570
  (
    .A(A[8]),
    .Y(n301)
  );


  sky130_fd_sc_hd__clkinv_1
  U1571
  (
    .A(n1643),
    .Y(n1605)
  );


  sky130_fd_sc_hd__xor2_1
  U1572
  (
    .A(n1623),
    .B(n872),
    .X(n1643)
  );


  sky130_fd_sc_hd__clkinv_1
  U1573
  (
    .A(n851),
    .Y(n872)
  );


  sky130_fd_sc_hd__nand2_1
  U1574
  (
    .A(A[7]),
    .B(n300),
    .Y(n1623)
  );


  sky130_fd_sc_hd__nand2_1
  U1575
  (
    .A(A[6]),
    .B(n300),
    .Y(n851)
  );


  sky130_fd_sc_hd__xnor2_1
  U1576
  (
    .A(n1627),
    .B(n1628),
    .Y(n1635)
  );


  sky130_fd_sc_hd__xnor2_1
  U1577
  (
    .A(n1145),
    .B(n1320),
    .Y(n1628)
  );


  sky130_fd_sc_hd__a221oi_1
  U1578
  (
    .A1(n1253),
    .A2(n1260),
    .B1(n1251),
    .B2(B[13]),
    .C1(n1645),
    .Y(n1320)
  );


  sky130_fd_sc_hd__o22ai_1
  U1579
  (
    .A1(n1154),
    .A2(n1385),
    .B1(n1262),
    .B2(n1351),
    .Y(n1645)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1580
  (
    .B1(n1646),
    .B2(n1647),
    .A1_N(n1648),
    .A2_N(n1322),
    .Y(n1627)
  );


  sky130_fd_sc_hd__nor2_1
  U1581
  (
    .A(n1647),
    .B(n1646),
    .Y(n1648)
  );


  sky130_fd_sc_hd__maj3_1
  U1582
  (
    .A(n1649),
    .B(n131),
    .C(n1650),
    .X(n1630)
  );


  sky130_fd_sc_hd__xor2_1
  U1583
  (
    .A(A[15]),
    .B(n442),
    .X(n1650)
  );


  sky130_fd_sc_hd__a221oi_1
  U1584
  (
    .A1(n1424),
    .A2(B[9]),
    .B1(n1393),
    .B2(n1152),
    .C1(n1651),
    .Y(n442)
  );


  sky130_fd_sc_hd__o22ai_1
  U1585
  (
    .A1(n1154),
    .A2(n1357),
    .B1(n1029),
    .B2(n1426),
    .Y(n1651)
  );


  sky130_fd_sc_hd__xor2_1
  U1586
  (
    .A(n1652),
    .B(n1653),
    .X(n1152)
  );


  sky130_fd_sc_hd__xor2_1
  U1587
  (
    .A(B[9]),
    .B(B[10]),
    .X(n1653)
  );


  sky130_fd_sc_hd__xnor2_1
  U1588
  (
    .A(n1654),
    .B(n1322),
    .Y(n131)
  );


  sky130_fd_sc_hd__xnor2_1
  U1589
  (
    .A(n1640),
    .B(n1641),
    .Y(n1322)
  );


  sky130_fd_sc_hd__xnor2_1
  U1590
  (
    .A(n834),
    .B(n1655),
    .Y(n1641)
  );


  sky130_fd_sc_hd__a221oi_1
  U1591
  (
    .A1(n1138),
    .A2(B[16]),
    .B1(n1164),
    .B2(B[15]),
    .C1(n1656),
    .Y(n1655)
  );


  sky130_fd_sc_hd__o22ai_1
  U1592
  (
    .A1(n1435),
    .A2(n1022),
    .B1(n1436),
    .B2(n1023),
    .Y(n1656)
  );


  sky130_fd_sc_hd__clkinv_1
  U1593
  (
    .A(n1137),
    .Y(n1022)
  );


  sky130_fd_sc_hd__nor3_1
  U1594
  (
    .A(n1657),
    .B(n1658),
    .C(n1659),
    .Y(n1137)
  );


  sky130_fd_sc_hd__nand3_1
  U1595
  (
    .A(A[9]),
    .B(n1660),
    .C(n1661),
    .Y(n1640)
  );


  sky130_fd_sc_hd__xnor2_1
  U1596
  (
    .A(n1647),
    .B(n1646),
    .Y(n1654)
  );


  sky130_fd_sc_hd__o22ai_1
  U1597
  (
    .A1(n1325),
    .A2(n1662),
    .B1(n1663),
    .B2(n1326),
    .Y(n1646)
  );


  sky130_fd_sc_hd__and2_0
  U1598
  (
    .A(n1662),
    .B(n1325),
    .X(n1663)
  );


  sky130_fd_sc_hd__xnor2_1
  U1599
  (
    .A(A[12]),
    .B(n1324),
    .Y(n1647)
  );


  sky130_fd_sc_hd__a221oi_1
  U1600
  (
    .A1(n1253),
    .A2(n1337),
    .B1(n1251),
    .B2(B[14]),
    .C1(n1664),
    .Y(n1324)
  );


  sky130_fd_sc_hd__o22ai_1
  U1601
  (
    .A1(n1262),
    .A2(n1385),
    .B1(n1185),
    .B2(n1351),
    .Y(n1664)
  );


  sky130_fd_sc_hd__maj3_1
  U1602
  (
    .A(n1665),
    .B(n127),
    .C(n1666),
    .X(n1649)
  );


  sky130_fd_sc_hd__xor2_1
  U1603
  (
    .A(A[15]),
    .B(n444),
    .X(n1666)
  );


  sky130_fd_sc_hd__a221oi_1
  U1604
  (
    .A1(n1393),
    .A2(n1187),
    .B1(n1391),
    .B2(B[12]),
    .C1(n1667),
    .Y(n444)
  );


  sky130_fd_sc_hd__o22ai_1
  U1605
  (
    .A1(n1029),
    .A2(n1457),
    .B1(n1154),
    .B2(n1426),
    .Y(n1667)
  );


  sky130_fd_sc_hd__xnor2_1
  U1606
  (
    .A(n1668),
    .B(n1669),
    .Y(n1187)
  );


  sky130_fd_sc_hd__xor2_1
  U1607
  (
    .A(B[11]),
    .B(B[10]),
    .X(n1669)
  );


  sky130_fd_sc_hd__xnor2_1
  U1608
  (
    .A(n1670),
    .B(n1326),
    .Y(n127)
  );


  sky130_fd_sc_hd__xnor2_1
  U1609
  (
    .A(n1661),
    .B(n1671),
    .Y(n1326)
  );


  sky130_fd_sc_hd__nor2b_1
  U1610
  (
    .B_N(n1660),
    .A(n834),
    .Y(n1671)
  );


  sky130_fd_sc_hd__xor2_1
  U1611
  (
    .A(n834),
    .B(n1672),
    .X(n1661)
  );


  sky130_fd_sc_hd__a222oi_1
  U1612
  (
    .A1(n1139),
    .A2(n1467),
    .B1(n1138),
    .B2(B[17]),
    .C1(n1164),
    .C2(B[16]),
    .Y(n1672)
  );


  sky130_fd_sc_hd__clkinv_1
  U1613
  (
    .A(n1178),
    .Y(n1164)
  );


  sky130_fd_sc_hd__clkinv_1
  U1614
  (
    .A(n1166),
    .Y(n1138)
  );


  sky130_fd_sc_hd__nand2b_1
  U1615
  (
    .A_N(n1659),
    .B(n1657),
    .Y(n1166)
  );


  sky130_fd_sc_hd__xor2_1
  U1616
  (
    .A(A[10]),
    .B(A[11]),
    .X(n1657)
  );


  sky130_fd_sc_hd__clkinv_1
  U1617
  (
    .A(n1023),
    .Y(n1139)
  );


  sky130_fd_sc_hd__xnor2_1
  U1618
  (
    .A(n1662),
    .B(n1325),
    .Y(n1670)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1619
  (
    .B1(n1673),
    .B2(n1674),
    .A1_N(n1675),
    .A2_N(n1676),
    .Y(n1325)
  );


  sky130_fd_sc_hd__xnor2_1
  U1620
  (
    .A(n1145),
    .B(n1328),
    .Y(n1662)
  );


  sky130_fd_sc_hd__a221oi_1
  U1621
  (
    .A1(n1253),
    .A2(n1559),
    .B1(n1251),
    .B2(B[15]),
    .C1(n1677),
    .Y(n1328)
  );


  sky130_fd_sc_hd__o22ai_1
  U1622
  (
    .A1(n1185),
    .A2(n1385),
    .B1(n1336),
    .B2(n1351),
    .Y(n1677)
  );


  sky130_fd_sc_hd__maj3_1
  U1623
  (
    .A(n1678),
    .B(n123),
    .C(n1679),
    .X(n1665)
  );


  sky130_fd_sc_hd__xor2_1
  U1624
  (
    .A(A[15]),
    .B(n446),
    .X(n1679)
  );


  sky130_fd_sc_hd__a221oi_1
  U1625
  (
    .A1(n1393),
    .A2(n1260),
    .B1(n1391),
    .B2(B[13]),
    .C1(n1680),
    .Y(n446)
  );


  sky130_fd_sc_hd__o22ai_1
  U1626
  (
    .A1(n1154),
    .A2(n1457),
    .B1(n1262),
    .B2(n1426),
    .Y(n1680)
  );


  sky130_fd_sc_hd__xor2_1
  U1627
  (
    .A(n1681),
    .B(n1682),
    .X(n1260)
  );


  sky130_fd_sc_hd__xor2_1
  U1628
  (
    .A(B[12]),
    .B(B[11]),
    .X(n1682)
  );


  sky130_fd_sc_hd__xnor2_1
  U1629
  (
    .A(n1675),
    .B(n1683),
    .Y(n123)
  );


  sky130_fd_sc_hd__xor2_1
  U1630
  (
    .A(n1673),
    .B(n1676),
    .X(n1683)
  );


  sky130_fd_sc_hd__clkinv_1
  U1631
  (
    .A(n1674),
    .Y(n1676)
  );


  sky130_fd_sc_hd__xor2_1
  U1632
  (
    .A(n1145),
    .B(n1684),
    .X(n1674)
  );


  sky130_fd_sc_hd__a221oi_1
  U1633
  (
    .A1(n1253),
    .A2(n1638),
    .B1(n1251),
    .B2(B[16]),
    .C1(n1685),
    .Y(n1684)
  );


  sky130_fd_sc_hd__o22ai_1
  U1634
  (
    .A1(n1336),
    .A2(n1385),
    .B1(n1369),
    .B2(n1351),
    .Y(n1685)
  );


  sky130_fd_sc_hd__nor2_1
  U1635
  (
    .A(n1686),
    .B(n1687),
    .Y(n1673)
  );


  sky130_fd_sc_hd__xor2_1
  U1636
  (
    .A(n1660),
    .B(n834),
    .X(n1675)
  );


  sky130_fd_sc_hd__xnor2_1
  U1637
  (
    .A(n834),
    .B(n1688),
    .Y(n1660)
  );


  sky130_fd_sc_hd__a21oi_1
  U1638
  (
    .A1(n1023),
    .A2(n1178),
    .B1(n1435),
    .Y(n1688)
  );


  sky130_fd_sc_hd__nand2_1
  U1639
  (
    .A(n1658),
    .B(n1659),
    .Y(n1178)
  );


  sky130_fd_sc_hd__nand2b_1
  U1640
  (
    .A_N(n1658),
    .B(n1659),
    .Y(n1023)
  );


  sky130_fd_sc_hd__xor2_1
  U1641
  (
    .A(A[11]),
    .B(A[12]),
    .X(n1659)
  );


  sky130_fd_sc_hd__xnor2_1
  U1642
  (
    .A(A[10]),
    .B(A[9]),
    .Y(n1658)
  );


  sky130_fd_sc_hd__clkinv_1
  U1643
  (
    .A(A[9]),
    .Y(n834)
  );


  sky130_fd_sc_hd__maj3_1
  U1644
  (
    .A(n1689),
    .B(n109),
    .C(n1690),
    .X(n1678)
  );


  sky130_fd_sc_hd__xor2_1
  U1645
  (
    .A(A[15]),
    .B(n448),
    .X(n1690)
  );


  sky130_fd_sc_hd__a221oi_1
  U1646
  (
    .A1(n1393),
    .A2(n1337),
    .B1(n1391),
    .B2(B[14]),
    .C1(n1691),
    .Y(n448)
  );


  sky130_fd_sc_hd__o22ai_1
  U1647
  (
    .A1(n1262),
    .A2(n1457),
    .B1(n1185),
    .B2(n1426),
    .Y(n1691)
  );


  sky130_fd_sc_hd__xor2_1
  U1648
  (
    .A(n1692),
    .B(n1693),
    .X(n1337)
  );


  sky130_fd_sc_hd__xor2_1
  U1649
  (
    .A(n1262),
    .B(B[13]),
    .X(n1692)
  );


  sky130_fd_sc_hd__xnor2_1
  U1650
  (
    .A(n1686),
    .B(n1687),
    .Y(n109)
  );


  sky130_fd_sc_hd__xnor2_1
  U1651
  (
    .A(n1145),
    .B(n1694),
    .Y(n1687)
  );


  sky130_fd_sc_hd__a221oi_1
  U1652
  (
    .A1(n1252),
    .A2(B[16]),
    .B1(n1349),
    .B2(B[15]),
    .C1(n1695),
    .Y(n1694)
  );


  sky130_fd_sc_hd__o22ai_1
  U1653
  (
    .A1(n1435),
    .A2(n1179),
    .B1(n1436),
    .B2(n1180),
    .Y(n1695)
  );


  sky130_fd_sc_hd__clkinv_1
  U1654
  (
    .A(n1251),
    .Y(n1179)
  );


  sky130_fd_sc_hd__nor3_1
  U1655
  (
    .A(n1696),
    .B(n1697),
    .C(n1698),
    .Y(n1251)
  );


  sky130_fd_sc_hd__nand3_1
  U1656
  (
    .A(A[12]),
    .B(n1699),
    .C(n1700),
    .Y(n1686)
  );


  sky130_fd_sc_hd__maj3_1
  U1657
  (
    .A(n107),
    .B(n105),
    .C(n1701),
    .X(n1689)
  );


  sky130_fd_sc_hd__xor2_1
  U1658
  (
    .A(A[15]),
    .B(n450),
    .X(n1701)
  );


  sky130_fd_sc_hd__a221oi_1
  U1659
  (
    .A1(n1393),
    .A2(n1559),
    .B1(n1391),
    .B2(B[15]),
    .C1(n1702),
    .Y(n450)
  );


  sky130_fd_sc_hd__o22ai_1
  U1660
  (
    .A1(n1185),
    .A2(n1457),
    .B1(n1336),
    .B2(n1426),
    .Y(n1702)
  );


  sky130_fd_sc_hd__xor2_1
  U1661
  (
    .A(n1703),
    .B(n1704),
    .X(n1559)
  );


  sky130_fd_sc_hd__xor2_1
  U1662
  (
    .A(B[14]),
    .B(B[13]),
    .X(n1704)
  );


  sky130_fd_sc_hd__xnor2_1
  U1663
  (
    .A(n1700),
    .B(n1705),
    .Y(n105)
  );


  sky130_fd_sc_hd__nor2b_1
  U1664
  (
    .B_N(n1699),
    .A(n1145),
    .Y(n1705)
  );


  sky130_fd_sc_hd__xor2_1
  U1665
  (
    .A(n1145),
    .B(n1706),
    .X(n1700)
  );


  sky130_fd_sc_hd__a222oi_1
  U1666
  (
    .A1(n1253),
    .A2(n1467),
    .B1(n1252),
    .B2(B[17]),
    .C1(n1349),
    .C2(B[16]),
    .Y(n1706)
  );


  sky130_fd_sc_hd__clkinv_1
  U1667
  (
    .A(n1385),
    .Y(n1349)
  );


  sky130_fd_sc_hd__clkinv_1
  U1668
  (
    .A(n1351),
    .Y(n1252)
  );


  sky130_fd_sc_hd__nand2_1
  U1669
  (
    .A(n1707),
    .B(n1696),
    .Y(n1351)
  );


  sky130_fd_sc_hd__xor2_1
  U1670
  (
    .A(A[13]),
    .B(A[14]),
    .X(n1696)
  );


  sky130_fd_sc_hd__a22oi_1
  U1671
  (
    .A1(n102),
    .A2(n101),
    .B1(n103),
    .B2(n101),
    .Y(n107)
  );


  sky130_fd_sc_hd__xor2_1
  U1672
  (
    .A(n1699),
    .B(A[12]),
    .X(n103)
  );


  sky130_fd_sc_hd__xnor2_1
  U1673
  (
    .A(n1145),
    .B(n1708),
    .Y(n1699)
  );


  sky130_fd_sc_hd__a21oi_1
  U1674
  (
    .A1(n1180),
    .A2(n1385),
    .B1(n1435),
    .Y(n1708)
  );


  sky130_fd_sc_hd__nand2_1
  U1675
  (
    .A(n1697),
    .B(n1698),
    .Y(n1385)
  );


  sky130_fd_sc_hd__clkinv_1
  U1676
  (
    .A(n1253),
    .Y(n1180)
  );


  sky130_fd_sc_hd__nor2_1
  U1677
  (
    .A(n1707),
    .B(n1697),
    .Y(n1253)
  );


  sky130_fd_sc_hd__xnor2_1
  U1678
  (
    .A(A[13]),
    .B(A[12]),
    .Y(n1697)
  );


  sky130_fd_sc_hd__clkinv_1
  U1679
  (
    .A(n1698),
    .Y(n1707)
  );


  sky130_fd_sc_hd__xor2_1
  U1680
  (
    .A(A[14]),
    .B(A[15]),
    .X(n1698)
  );


  sky130_fd_sc_hd__clkinv_1
  U1681
  (
    .A(A[12]),
    .Y(n1145)
  );


  sky130_fd_sc_hd__xnor2_1
  U1682
  (
    .A(A[15]),
    .B(n1709),
    .Y(n101)
  );


  sky130_fd_sc_hd__a221oi_1
  U1683
  (
    .A1(n1393),
    .A2(n1638),
    .B1(n1391),
    .B2(B[16]),
    .C1(n1710),
    .Y(n1709)
  );


  sky130_fd_sc_hd__o22ai_1
  U1684
  (
    .A1(n1336),
    .A2(n1457),
    .B1(n1369),
    .B2(n1426),
    .Y(n1710)
  );


  sky130_fd_sc_hd__clkinv_1
  U1685
  (
    .A(n1403),
    .Y(n1638)
  );


  sky130_fd_sc_hd__xor2_1
  U1686
  (
    .A(n1711),
    .B(n1712),
    .X(n1403)
  );


  sky130_fd_sc_hd__xor2_1
  U1687
  (
    .A(n1369),
    .B(B[14]),
    .X(n1711)
  );


  sky130_fd_sc_hd__nor2_1
  U1688
  (
    .A(n98),
    .B(n99),
    .Y(n102)
  );


  sky130_fd_sc_hd__xnor2_1
  U1689
  (
    .A(n97),
    .B(n1713),
    .Y(n99)
  );


  sky130_fd_sc_hd__a221oi_1
  U1690
  (
    .A1(n1392),
    .A2(B[16]),
    .B1(n1424),
    .B2(B[15]),
    .C1(n1714),
    .Y(n1713)
  );


  sky130_fd_sc_hd__o22ai_1
  U1691
  (
    .A1(n1435),
    .A2(n1357),
    .B1(n1436),
    .B2(n1358),
    .Y(n1714)
  );


  sky130_fd_sc_hd__xor2_1
  U1692
  (
    .A(n1715),
    .B(n1716),
    .X(n1436)
  );


  sky130_fd_sc_hd__xor2_1
  U1693
  (
    .A(B[16]),
    .B(B[15]),
    .X(n1716)
  );


  sky130_fd_sc_hd__clkinv_1
  U1694
  (
    .A(n1391),
    .Y(n1357)
  );


  sky130_fd_sc_hd__nor3b_1
  U1695
  (
    .C_N(n1717),
    .A(A[16]),
    .B(A[17]),
    .Y(n1391)
  );


  sky130_fd_sc_hd__nand3_1
  U1696
  (
    .A(A[15]),
    .B(n94),
    .C(n95),
    .Y(n98)
  );


  sky130_fd_sc_hd__xor2_1
  U1697
  (
    .A(n97),
    .B(n1718),
    .X(n95)
  );


  sky130_fd_sc_hd__a222oi_1
  U1698
  (
    .A1(n1393),
    .A2(n1467),
    .B1(n1392),
    .B2(B[17]),
    .C1(n1424),
    .C2(B[16]),
    .Y(n1718)
  );


  sky130_fd_sc_hd__clkinv_1
  U1699
  (
    .A(n1426),
    .Y(n1392)
  );


  sky130_fd_sc_hd__nand2_1
  U1700
  (
    .A(A[16]),
    .B(n1719),
    .Y(n1426)
  );


  sky130_fd_sc_hd__xor2_1
  U1701
  (
    .A(B[17]),
    .B(B[16]),
    .X(n1467)
  );


  sky130_fd_sc_hd__clkinv_1
  U1702
  (
    .A(n1358),
    .Y(n1393)
  );


  sky130_fd_sc_hd__xnor2_1
  U1703
  (
    .A(n97),
    .B(n1720),
    .Y(n94)
  );


  sky130_fd_sc_hd__a21oi_1
  U1704
  (
    .A1(n1358),
    .A2(n1457),
    .B1(n1435),
    .Y(n1720)
  );


  sky130_fd_sc_hd__clkinv_1
  U1705
  (
    .A(B[17]),
    .Y(n1435)
  );


  sky130_fd_sc_hd__clkinv_1
  U1706
  (
    .A(n1424),
    .Y(n1457)
  );


  sky130_fd_sc_hd__nor2_1
  U1707
  (
    .A(n1717),
    .B(n1719),
    .Y(n1424)
  );


  sky130_fd_sc_hd__clkinv_1
  U1708
  (
    .A(A[17]),
    .Y(n1719)
  );


  sky130_fd_sc_hd__nand2_1
  U1709
  (
    .A(A[17]),
    .B(n1717),
    .Y(n1358)
  );


  sky130_fd_sc_hd__xor2_1
  U1710
  (
    .A(A[16]),
    .B(A[15]),
    .X(n1717)
  );


  sky130_fd_sc_hd__clkinv_1
  U1711
  (
    .A(A[15]),
    .Y(n97)
  );


  sky130_fd_sc_hd__maj3_1
  U1712
  (
    .A(n754),
    .B(n755),
    .C(n236),
    .X(n742)
  );


  sky130_fd_sc_hd__nor2_1
  U1713
  (
    .A(n786),
    .B(n739),
    .Y(n236)
  );


  sky130_fd_sc_hd__nand2_1
  U1714
  (
    .A(n740),
    .B(n768),
    .Y(n755)
  );


  sky130_fd_sc_hd__clkinv_1
  U1715
  (
    .A(n788),
    .Y(n768)
  );


  sky130_fd_sc_hd__clkinv_1
  U1716
  (
    .A(n739),
    .Y(n740)
  );


  sky130_fd_sc_hd__xor2_1
  U1717
  (
    .A(n739),
    .B(n1721),
    .X(n754)
  );


  sky130_fd_sc_hd__o22ai_1
  U1718
  (
    .A1(n810),
    .A2(n787),
    .B1(n1370),
    .B2(n813),
    .Y(n1721)
  );


  sky130_fd_sc_hd__nand2_1
  U1719
  (
    .A(n741),
    .B(n1394),
    .Y(n813)
  );


  sky130_fd_sc_hd__o22ai_1
  U1720
  (
    .A1(n1427),
    .A2(n810),
    .B1(n1722),
    .B2(n788),
    .Y(n1394)
  );


  sky130_fd_sc_hd__nor2b_1
  U1721
  (
    .B_N(n1427),
    .A(n741),
    .Y(n1722)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1722
  (
    .B1(n1458),
    .B2(n1460),
    .A1_N(n1723),
    .A2_N(n788),
    .Y(n1427)
  );


  sky130_fd_sc_hd__nand2_1
  U1723
  (
    .A(B[1]),
    .B(n300),
    .Y(n788)
  );


  sky130_fd_sc_hd__nor2_1
  U1724
  (
    .A(n1460),
    .B(n1458),
    .Y(n1723)
  );


  sky130_fd_sc_hd__clkinv_1
  U1725
  (
    .A(n786),
    .Y(n1460)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1726
  (
    .B1(n1724),
    .B2(n786),
    .A1_N(n1490),
    .A2_N(n807),
    .Y(n1458)
  );


  sky130_fd_sc_hd__nand2_1
  U1727
  (
    .A(B[2]),
    .B(n300),
    .Y(n786)
  );


  sky130_fd_sc_hd__nor2_1
  U1728
  (
    .A(n807),
    .B(n1490),
    .Y(n1724)
  );


  sky130_fd_sc_hd__o22ai_1
  U1729
  (
    .A1(n1725),
    .A2(n815),
    .B1(n1726),
    .B2(n781),
    .Y(n1490)
  );


  sky130_fd_sc_hd__nor2_1
  U1730
  (
    .A(n1519),
    .B(n1517),
    .Y(n1726)
  );


  sky130_fd_sc_hd__clkinv_1
  U1731
  (
    .A(n815),
    .Y(n1519)
  );


  sky130_fd_sc_hd__clkinv_1
  U1732
  (
    .A(n1517),
    .Y(n1725)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1733
  (
    .B1(n1727),
    .B2(n815),
    .A1_N(n1544),
    .A2_N(n853),
    .Y(n1517)
  );


  sky130_fd_sc_hd__nand2_1
  U1734
  (
    .A(B[4]),
    .B(n300),
    .Y(n815)
  );


  sky130_fd_sc_hd__nor2_1
  U1735
  (
    .A(n853),
    .B(n1544),
    .Y(n1727)
  );


  sky130_fd_sc_hd__o22ai_1
  U1736
  (
    .A1(n1571),
    .A2(n873),
    .B1(n1728),
    .B2(n876),
    .Y(n1544)
  );


  sky130_fd_sc_hd__nor2b_1
  U1737
  (
    .B_N(n1571),
    .A(n908),
    .Y(n1728)
  );


  sky130_fd_sc_hd__clkinv_1
  U1738
  (
    .A(n873),
    .Y(n908)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1739
  (
    .B1(n1592),
    .B2(n905),
    .A1_N(n1729),
    .A2_N(n873),
    .Y(n1571)
  );


  sky130_fd_sc_hd__nand2_1
  U1740
  (
    .A(B[6]),
    .B(n300),
    .Y(n873)
  );


  sky130_fd_sc_hd__nor2_1
  U1741
  (
    .A(n905),
    .B(n1592),
    .Y(n1729)
  );


  sky130_fd_sc_hd__clkinv_1
  U1742
  (
    .A(n1037),
    .Y(n905)
  );


  sky130_fd_sc_hd__o22ai_1
  U1743
  (
    .A1(n1730),
    .A2(n970),
    .B1(n1731),
    .B2(n1037),
    .Y(n1592)
  );


  sky130_fd_sc_hd__nand2_1
  U1744
  (
    .A(B[7]),
    .B(n300),
    .Y(n1037)
  );


  sky130_fd_sc_hd__nor2_1
  U1745
  (
    .A(n1732),
    .B(n1616),
    .Y(n1731)
  );


  sky130_fd_sc_hd__clkinv_1
  U1746
  (
    .A(n1616),
    .Y(n1730)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1747
  (
    .B1(n1733),
    .B2(n993),
    .A1_N(n1633),
    .A2_N(n1732),
    .Y(n1616)
  );


  sky130_fd_sc_hd__nor2_1
  U1748
  (
    .A(n1732),
    .B(n1633),
    .Y(n1733)
  );


  sky130_fd_sc_hd__o2bb2ai_1
  U1749
  (
    .B1(n1734),
    .B2(n993),
    .A1_N(n1652),
    .A2_N(B[10]),
    .Y(n1633)
  );


  sky130_fd_sc_hd__clkinv_1
  U1750
  (
    .A(B[9]),
    .Y(n993)
  );


  sky130_fd_sc_hd__nor2_1
  U1751
  (
    .A(B[10]),
    .B(n1652),
    .Y(n1734)
  );


  sky130_fd_sc_hd__o22ai_1
  U1752
  (
    .A1(n1668),
    .A2(n1029),
    .B1(n1735),
    .B2(n1154),
    .Y(n1652)
  );


  sky130_fd_sc_hd__clkinv_1
  U1753
  (
    .A(B[11]),
    .Y(n1154)
  );


  sky130_fd_sc_hd__nor2b_1
  U1754
  (
    .B_N(n1668),
    .A(B[10]),
    .Y(n1735)
  );


  sky130_fd_sc_hd__clkinv_1
  U1755
  (
    .A(B[10]),
    .Y(n1029)
  );


  sky130_fd_sc_hd__a21boi_0
  U1756
  (
    .A1(n1681),
    .A2(B[11]),
    .B1_N(n1736),
    .Y(n1668)
  );


  sky130_fd_sc_hd__o21ai_0
  U1757
  (
    .A1(B[11]),
    .A2(n1681),
    .B1(B[12]),
    .Y(n1736)
  );


  sky130_fd_sc_hd__o22ai_1
  U1758
  (
    .A1(n1693),
    .A2(n1262),
    .B1(n1737),
    .B2(n1185),
    .Y(n1681)
  );


  sky130_fd_sc_hd__clkinv_1
  U1759
  (
    .A(B[13]),
    .Y(n1185)
  );


  sky130_fd_sc_hd__nor2b_1
  U1760
  (
    .B_N(n1693),
    .A(B[12]),
    .Y(n1737)
  );


  sky130_fd_sc_hd__clkinv_1
  U1761
  (
    .A(B[12]),
    .Y(n1262)
  );


  sky130_fd_sc_hd__a2bb2oi_1
  U1762
  (
    .B1(n1703),
    .B2(B[13]),
    .A1_N(n1738),
    .A2_N(n1336),
    .Y(n1693)
  );


  sky130_fd_sc_hd__clkinv_1
  U1763
  (
    .A(B[14]),
    .Y(n1336)
  );


  sky130_fd_sc_hd__nor2_1
  U1764
  (
    .A(B[13]),
    .B(n1703),
    .Y(n1738)
  );


  sky130_fd_sc_hd__maj3_1
  U1765
  (
    .A(n1712),
    .B(B[15]),
    .C(B[14]),
    .X(n1703)
  );


  sky130_fd_sc_hd__a21oi_1
  U1766
  (
    .A1(n1715),
    .A2(n1369),
    .B1(n1402),
    .Y(n1712)
  );


  sky130_fd_sc_hd__clkinv_1
  U1767
  (
    .A(B[16]),
    .Y(n1402)
  );


  sky130_fd_sc_hd__clkinv_1
  U1768
  (
    .A(B[15]),
    .Y(n1369)
  );


  sky130_fd_sc_hd__nand2_1
  U1769
  (
    .A(B[17]),
    .B(B[16]),
    .Y(n1715)
  );


  sky130_fd_sc_hd__clkinv_1
  U1770
  (
    .A(n970),
    .Y(n1732)
  );


  sky130_fd_sc_hd__nand2_1
  U1771
  (
    .A(B[8]),
    .B(n300),
    .Y(n970)
  );


  sky130_fd_sc_hd__clkinv_1
  U1772
  (
    .A(n876),
    .Y(n853)
  );


  sky130_fd_sc_hd__nand2_1
  U1773
  (
    .A(B[5]),
    .B(n300),
    .Y(n876)
  );


  sky130_fd_sc_hd__clkinv_1
  U1774
  (
    .A(n781),
    .Y(n807)
  );


  sky130_fd_sc_hd__nand2_1
  U1775
  (
    .A(B[3]),
    .B(n300),
    .Y(n781)
  );


  sky130_fd_sc_hd__clkinv_1
  U1776
  (
    .A(n810),
    .Y(n741)
  );


  sky130_fd_sc_hd__clkinv_1
  U1777
  (
    .A(n771),
    .Y(n1370)
  );


  sky130_fd_sc_hd__nor2b_1
  U1778
  (
    .B_N(n1501),
    .A(n1468),
    .Y(n771)
  );


  sky130_fd_sc_hd__nand3b_1
  U1779
  (
    .A_N(n1469),
    .B(n1501),
    .C(n1468),
    .Y(n787)
  );


  sky130_fd_sc_hd__xor2_1
  U1780
  (
    .A(n751),
    .B(n1739),
    .X(n1468)
  );


  sky130_fd_sc_hd__nand2_1
  U1781
  (
    .A(A[3]),
    .B(n300),
    .Y(n751)
  );


  sky130_fd_sc_hd__xnor2_1
  U1782
  (
    .A(n739),
    .B(n1740),
    .Y(n1501)
  );


  sky130_fd_sc_hd__xor2_1
  U1783
  (
    .A(n1740),
    .B(n1739),
    .X(n1469)
  );


  sky130_fd_sc_hd__nor2_1
  U1784
  (
    .A(n733),
    .B(MODE_0_0),
    .Y(n1739)
  );


  sky130_fd_sc_hd__clkinv_1
  U1785
  (
    .A(A[2]),
    .Y(n733)
  );


  sky130_fd_sc_hd__nor2_1
  U1786
  (
    .A(n498),
    .B(MODE_0_0),
    .Y(n1740)
  );


  sky130_fd_sc_hd__clkinv_1
  U1787
  (
    .A(A[1]),
    .Y(n498)
  );


  sky130_fd_sc_hd__nand2_1
  U1788
  (
    .A(B[0]),
    .B(n300),
    .Y(n810)
  );


  sky130_fd_sc_hd__nand2_1
  U1789
  (
    .A(A[0]),
    .B(n300),
    .Y(n739)
  );


  sky130_fd_sc_hd__clkinv_1
  U1790
  (
    .A(MODE_0_0),
    .Y(n300)
  );


endmodule

