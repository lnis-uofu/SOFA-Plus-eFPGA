

module direct_interc
(
  input [0:0] in,
  output [0:0] out
);

  wire [0:0] in;
  wire [0:0] out;
  assign out[0] = in[0];

endmodule

