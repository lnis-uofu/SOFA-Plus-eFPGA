

module sb_0__3_
( config_enable, pReset, chany_top_in, top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_, chany_bottom_in, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, ccff_head, chany_top_out, chanx_right_out, chany_bottom_out, ccff_tail, pReset_E_in, pReset_S_out, config_enable_E_in, config_enable_S_out, prog_clk, prog_clk_0_E_in ); 
  input [0:0] config_enable;
  input [0:0] pReset;
  input [0:19] chany_top_in;
  input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
  input [0:19] chanx_right_in;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_;
  input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_;
  input [0:19] chany_bottom_in;
  input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
  input [0:0] ccff_head;
  output [0:19] chany_top_out;
  output [0:19] chanx_right_out;
  output [0:19] chany_bottom_out;
  output [0:0] ccff_tail;
  input pReset_E_in;
  output pReset_S_out;
  input config_enable_E_in;
  output config_enable_S_out;
  input prog_clk;
  input prog_clk_0_E_in;

  wire [0:1] mux_tree_tapbuf_size2_0_sram;
  wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
  wire [0:1] mux_tree_tapbuf_size2_1_sram;
  wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
  wire [0:1] mux_tree_tapbuf_size2_2_sram;
  wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
  wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
  wire [0:1] mux_tree_tapbuf_size3_0_sram;
  wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_1_sram;
  wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_2_sram;
  wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_3_sram;
  wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_4_sram;
  wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_5_sram;
  wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_6_sram;
  wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
  wire [0:1] mux_tree_tapbuf_size3_7_sram;
  wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
  wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
  wire [0:2] mux_tree_tapbuf_size4_0_sram;
  wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
  wire [0:2] mux_tree_tapbuf_size4_1_sram;
  wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
  wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
  wire [0:2] mux_tree_tapbuf_size5_0_sram;
  wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_1_sram;
  wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_2_sram;
  wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_3_sram;
  wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_4_sram;
  wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_5_sram;
  wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_6_sram;
  wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_7_sram;
  wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_8_sram;
  wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
  wire [0:2] mux_tree_tapbuf_size5_9_sram;
  wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
  wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
  wire [0:2] mux_tree_tapbuf_size6_0_sram;
  wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
  wire [0:2] mux_tree_tapbuf_size6_1_sram;
  wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
  wire [0:2] mux_tree_tapbuf_size6_2_sram;
  wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
  wire [0:2] mux_tree_tapbuf_size6_3_sram;
  wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
  wire [0:2] mux_tree_tapbuf_size6_4_sram;
  wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
  wire [0:2] mux_tree_tapbuf_size6_5_sram;
  wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
  wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
  wire [0:3] mux_tree_tapbuf_size8_0_sram;
  wire [0:3] mux_tree_tapbuf_size8_0_sram_inv;
  wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail;
  wire [0:3] mux_tree_tapbuf_size9_0_sram;
  wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
  wire [0:3] mux_tree_tapbuf_size9_1_sram;
  wire [0:3] mux_tree_tapbuf_size9_1_sram_inv;
  wire [0:3] mux_tree_tapbuf_size9_2_sram;
  wire [0:3] mux_tree_tapbuf_size9_2_sram_inv;
  wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail;
  wire [0:0] mux_tree_tapbuf_size9_mem_2_ccff_tail;
  wire prog_clk_0;
  assign chany_bottom_out[3] = chany_top_in[2];
  assign chany_bottom_out[5] = chany_top_in[4];
  assign chany_bottom_out[6] = chany_top_in[5];
  assign chany_bottom_out[7] = chany_top_in[6];
  assign chany_bottom_out[9] = chany_top_in[8];
  assign chany_bottom_out[10] = chany_top_in[9];
  assign chany_bottom_out[11] = chany_top_in[10];
  assign chany_bottom_out[13] = chany_top_in[12];
  assign chany_bottom_out[14] = chany_top_in[13];
  assign chany_bottom_out[15] = chany_top_in[14];
  assign chany_bottom_out[17] = chany_top_in[16];
  assign chany_bottom_out[18] = chany_top_in[17];
  assign chany_bottom_out[19] = chany_top_in[18];
  assign chanx_right_out[19] = right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_[0];
  assign chany_top_out[3] = chany_bottom_in[2];
  assign chany_top_out[5] = chany_bottom_in[4];
  assign chany_top_out[6] = chany_bottom_in[5];
  assign chany_top_out[7] = chany_bottom_in[6];
  assign chany_top_out[9] = chany_bottom_in[8];
  assign chany_top_out[10] = chany_bottom_in[9];
  assign chany_top_out[11] = chany_bottom_in[10];
  assign chany_top_out[13] = chany_bottom_in[12];
  assign chany_top_out[14] = chany_bottom_in[13];
  assign chany_top_out[15] = chany_bottom_in[14];
  assign chany_top_out[17] = chany_bottom_in[16];
  assign chany_top_out[18] = chany_bottom_in[17];
  assign chany_top_out[19] = chany_bottom_in[18];
  assign prog_clk = prog_clk_0;

  mux_tree_tapbuf_size6
  mux_top_track_0
  (
    .in({ top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[1], chanx_right_in[8], chanx_right_in[15], chany_bottom_in[2], chany_bottom_in[12] }),
    .sram(mux_tree_tapbuf_size6_0_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
    .out(chany_top_out[0])
  );


  mux_tree_tapbuf_size6
  mux_top_track_4
  (
    .in({ top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[3], chanx_right_in[10], chanx_right_in[17], chany_bottom_in[5], chany_bottom_in[14] }),
    .sram(mux_tree_tapbuf_size6_1_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
    .out(chany_top_out[2])
  );


  mux_tree_tapbuf_size6
  mux_top_track_8
  (
    .in({ top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[4], chanx_right_in[11], chanx_right_in[18], chany_bottom_in[6], chany_bottom_in[16] }),
    .sram(mux_tree_tapbuf_size6_2_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
    .out(chany_top_out[4])
  );


  mux_tree_tapbuf_size6
  mux_bottom_track_1
  (
    .in({ chany_top_in[2], chany_top_in[12], chanx_right_in[5], chanx_right_in[12], chanx_right_in[19], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ }),
    .sram(mux_tree_tapbuf_size6_3_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
    .out(chany_bottom_out[0])
  );


  mux_tree_tapbuf_size6
  mux_bottom_track_5
  (
    .in({ chany_top_in[5], chany_top_in[14], chanx_right_in[3], chanx_right_in[10], chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ }),
    .sram(mux_tree_tapbuf_size6_4_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
    .out(chany_bottom_out[2])
  );


  mux_tree_tapbuf_size6
  mux_bottom_track_9
  (
    .in({ chany_top_in[6], chany_top_in[16], chanx_right_in[2], chanx_right_in[9], chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ }),
    .sram(mux_tree_tapbuf_size6_5_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
    .out(chany_bottom_out[4])
  );


  mux_tree_tapbuf_size6_mem
  mem_top_track_0
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(ccff_head),
    .ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2])
  );


  mux_tree_tapbuf_size6_mem
  mem_top_track_4
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2])
  );


  mux_tree_tapbuf_size6_mem
  mem_top_track_8
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2])
  );


  mux_tree_tapbuf_size6_mem
  mem_bottom_track_1
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2])
  );


  mux_tree_tapbuf_size6_mem
  mem_bottom_track_5
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2])
  );


  mux_tree_tapbuf_size6_mem
  mem_bottom_track_9
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
    .mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5
  mux_top_track_2
  (
    .in({ chanx_right_in[2], chanx_right_in[9], chanx_right_in[16], chany_bottom_in[4], chany_bottom_in[13] }),
    .sram(mux_tree_tapbuf_size5_0_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
    .out(chany_top_out[1])
  );


  mux_tree_tapbuf_size5
  mux_top_track_16
  (
    .in({ chanx_right_in[5], chanx_right_in[12], chanx_right_in[19], chany_bottom_in[8], chany_bottom_in[17] }),
    .sram(mux_tree_tapbuf_size5_1_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
    .out(chany_top_out[8])
  );


  mux_tree_tapbuf_size5
  mux_right_track_8
  (
    .in({ chany_top_in[7:8], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_, chany_bottom_in[8] }),
    .sram(mux_tree_tapbuf_size5_2_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
    .out(chanx_right_out[4])
  );


  mux_tree_tapbuf_size5
  mux_right_track_10
  (
    .in({ chany_top_in[9], chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_, chany_bottom_in[9] }),
    .sram(mux_tree_tapbuf_size5_3_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
    .out(chanx_right_out[5])
  );


  mux_tree_tapbuf_size5
  mux_right_track_12
  (
    .in({ chany_top_in[10], chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_, chany_bottom_in[10] }),
    .sram(mux_tree_tapbuf_size5_4_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
    .out(chanx_right_out[6])
  );


  mux_tree_tapbuf_size5
  mux_right_track_14
  (
    .in({ chany_top_in[12], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_, chany_bottom_in[12] }),
    .sram(mux_tree_tapbuf_size5_5_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
    .out(chanx_right_out[7])
  );


  mux_tree_tapbuf_size5
  mux_right_track_24
  (
    .in({ chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_, chany_bottom_in[18:19] }),
    .sram(mux_tree_tapbuf_size5_6_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
    .out(chanx_right_out[12])
  );


  mux_tree_tapbuf_size5
  mux_bottom_track_3
  (
    .in({ chany_top_in[4], chany_top_in[13], chanx_right_in[4], chanx_right_in[11], chanx_right_in[18] }),
    .sram(mux_tree_tapbuf_size5_7_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
    .out(chany_bottom_out[1])
  );


  mux_tree_tapbuf_size5
  mux_bottom_track_17
  (
    .in({ chany_top_in[8], chany_top_in[17], chanx_right_in[1], chanx_right_in[8], chanx_right_in[15] }),
    .sram(mux_tree_tapbuf_size5_8_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
    .out(chany_bottom_out[8])
  );


  mux_tree_tapbuf_size5
  mux_bottom_track_25
  (
    .in({ chany_top_in[9], chany_top_in[18], chanx_right_in[0], chanx_right_in[7], chanx_right_in[14] }),
    .sram(mux_tree_tapbuf_size5_9_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
    .out(chany_bottom_out[12])
  );


  mux_tree_tapbuf_size5_mem
  mem_top_track_2
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_top_track_16
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_right_track_8
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size9_mem_2_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_right_track_10
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_right_track_12
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_right_track_14
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_right_track_24
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_bottom_track_3
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_bottom_track_17
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2])
  );


  mux_tree_tapbuf_size5_mem
  mem_bottom_track_25
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
    .mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2])
  );


  mux_tree_tapbuf_size4
  mux_top_track_24
  (
    .in({ chanx_right_in[6], chanx_right_in[13], chany_bottom_in[9], chany_bottom_in[18] }),
    .sram(mux_tree_tapbuf_size4_0_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
    .out(chany_top_out[12])
  );


  mux_tree_tapbuf_size4
  mux_top_track_32
  (
    .in({ chanx_right_in[0], chanx_right_in[7], chanx_right_in[14], chany_bottom_in[10] }),
    .sram(mux_tree_tapbuf_size4_1_sram[0:2]),
    .sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
    .out(chany_top_out[16])
  );


  mux_tree_tapbuf_size4_mem
  mem_top_track_24
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2])
  );


  mux_tree_tapbuf_size4_mem
  mem_top_track_32
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
    .mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2])
  );


  mux_tree_tapbuf_size8
  mux_right_track_0
  (
    .in({ chany_top_in[2], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_, chany_bottom_in[2] }),
    .sram(mux_tree_tapbuf_size8_0_sram[0:3]),
    .sram_inv(mux_tree_tapbuf_size8_0_sram_inv[0:3]),
    .out(chanx_right_out[0])
  );


  mux_tree_tapbuf_size8_mem
  mem_right_track_0
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size8_0_sram[0:3]),
    .mem_outb(mux_tree_tapbuf_size8_0_sram_inv[0:3])
  );


  mux_tree_tapbuf_size9
  mux_right_track_2
  (
    .in({ chany_top_in[0], chany_top_in[4], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_, chany_bottom_in[4] }),
    .sram(mux_tree_tapbuf_size9_0_sram[0:3]),
    .sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
    .out(chanx_right_out[1])
  );


  mux_tree_tapbuf_size9
  mux_right_track_4
  (
    .in({ chany_top_in[1], chany_top_in[5], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_, chany_bottom_in[5] }),
    .sram(mux_tree_tapbuf_size9_1_sram[0:3]),
    .sram_inv(mux_tree_tapbuf_size9_1_sram_inv[0:3]),
    .out(chanx_right_out[2])
  );


  mux_tree_tapbuf_size9
  mux_right_track_6
  (
    .in({ chany_top_in[3], chany_top_in[6], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_, chany_bottom_in[6] }),
    .sram(mux_tree_tapbuf_size9_2_sram[0:3]),
    .sram_inv(mux_tree_tapbuf_size9_2_sram_inv[0:3]),
    .out(chanx_right_out[3])
  );


  mux_tree_tapbuf_size9_mem
  mem_right_track_2
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
    .mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3])
  );


  mux_tree_tapbuf_size9_mem
  mem_right_track_4
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size9_1_sram[0:3]),
    .mem_outb(mux_tree_tapbuf_size9_1_sram_inv[0:3])
  );


  mux_tree_tapbuf_size9_mem
  mem_right_track_6
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size9_mem_2_ccff_tail),
    .mem_out(mux_tree_tapbuf_size9_2_sram[0:3]),
    .mem_outb(mux_tree_tapbuf_size9_2_sram_inv[0:3])
  );


  mux_tree_tapbuf_size3
  mux_right_track_16
  (
    .in({ chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_, chany_bottom_in[13] }),
    .sram(mux_tree_tapbuf_size3_0_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
    .out(chanx_right_out[8])
  );


  mux_tree_tapbuf_size3
  mux_right_track_18
  (
    .in({ chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_, chany_bottom_in[14] }),
    .sram(mux_tree_tapbuf_size3_1_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
    .out(chanx_right_out[9])
  );


  mux_tree_tapbuf_size3
  mux_right_track_20
  (
    .in({ chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_, chany_bottom_in[16] }),
    .sram(mux_tree_tapbuf_size3_2_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
    .out(chanx_right_out[10])
  );


  mux_tree_tapbuf_size3
  mux_right_track_22
  (
    .in({ chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_7_, chany_bottom_in[17] }),
    .sram(mux_tree_tapbuf_size3_3_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
    .out(chanx_right_out[11])
  );


  mux_tree_tapbuf_size3
  mux_right_track_26
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_9_, chany_bottom_in[15] }),
    .sram(mux_tree_tapbuf_size3_4_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
    .out(chanx_right_out[13])
  );


  mux_tree_tapbuf_size3
  mux_right_track_28
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_10_, chany_bottom_in[11] }),
    .sram(mux_tree_tapbuf_size3_5_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
    .out(chanx_right_out[14])
  );


  mux_tree_tapbuf_size3
  mux_right_track_30
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_11_, chany_bottom_in[7] }),
    .sram(mux_tree_tapbuf_size3_6_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
    .out(chanx_right_out[15])
  );


  mux_tree_tapbuf_size3
  mux_bottom_track_33
  (
    .in({ chany_top_in[10], chanx_right_in[6], chanx_right_in[13] }),
    .sram(mux_tree_tapbuf_size3_7_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
    .out(chany_bottom_out[16])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_16
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_18
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_20
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_22
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_26
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_28
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_right_track_30
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1])
  );


  mux_tree_tapbuf_size3_mem
  mem_bottom_track_33
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
    .ccff_tail(ccff_tail),
    .mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1])
  );


  mux_tree_tapbuf_size2
  mux_right_track_32
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_4_, chany_bottom_in[3] }),
    .sram(mux_tree_tapbuf_size2_0_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
    .out(chanx_right_out[16])
  );


  mux_tree_tapbuf_size2
  mux_right_track_34
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_5_, chany_bottom_in[1] }),
    .sram(mux_tree_tapbuf_size2_1_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
    .out(chanx_right_out[17])
  );


  mux_tree_tapbuf_size2
  mux_right_track_36
  (
    .in({ right_bottom_grid_top_width_0_height_0_subtile_0__pin_out_6_, chany_bottom_in[0] }),
    .sram(mux_tree_tapbuf_size2_2_sram[0:1]),
    .sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
    .out(chanx_right_out[18])
  );


  mux_tree_tapbuf_size2_mem
  mem_right_track_32
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
    .mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1])
  );


  mux_tree_tapbuf_size2_mem
  mem_right_track_34
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
    .mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1])
  );


  mux_tree_tapbuf_size2_mem
  mem_right_track_36
  (
    .config_enable(config_enable),
    .pReset(pReset),
    .prog_clk(prog_clk),
    .ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
    .ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
    .mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
    .mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1])
  );


  BUF_X8
  pReset_FTB00
  (
    .A(pReset_E_in),
    .Y(pReset)
  );


  BUFCLK_X4
  pReset_S_FTB01
  (
    .A(pReset_E_in),
    .Y(pReset_S_out)
  );


  BUF_X8
  config_enable_FTB00
  (
    .A(config_enable_E_in),
    .Y(config_enable)
  );


  BUFCLK_X4
  config_enable_S_FTB01
  (
    .A(config_enable_E_in),
    .Y(config_enable_S_out)
  );


  BUF_X8
  prog_clk_0_FTB00
  (
    .A(prog_clk_0_E_in),
    .Y(prog_clk_0)
  );


endmodule

