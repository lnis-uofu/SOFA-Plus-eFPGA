//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Fabric Netlist Summary
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ------ Include defines: preproc flags -----
`include "./SRC/fpga_defines.v"

// ------ Include user-defined netlists -----
`include "./inv/sky130_fd_sc_hd__inv_1.v"
`include "./SRC/CustomModules/sky130_fd_sc_hd_wrapper.v"
`include "./SRC/CustomModules/sofa_plus_dff.v"
`include "./SRC/CustomModules/frac_lut4_arith.v"
`include "./SRC/CustomModules/sofa_plus_ccff.v"
`include "./SRC/CustomModules/sofa_plus_io.v"
`include "./RTL/frac_mult_18x18.v"
// ------ Include primitive module netlists -----
`include "./SRC/sub_module/inv_buf_passgate.v"
`include "./SRC/sub_module/arch_encoder.v"
`include "./SRC/sub_module/local_encoder.v"
`include "./SRC/sub_module/mux_primitives.v"
`include "./SRC/sub_module/muxes.v"
`include "./SRC/sub_module/luts.v"
`include "./SRC/sub_module/wires.v"
`include "./SRC/sub_module/memories.v"
`include "./SRC/sub_module/CBxFeedthrough.v"
`include "./SRC/sub_module/CByFeedthrough.v"
`include "./SRC/sub_module/CLBFeedthrough.v"

// ------ Include logic block netlists -----
`include "./SRC/lb/logical_tile_io_mode_physical__iopad.v"
`include "./SRC/lb/logical_tile_io_mode_io_.v"
`include "./SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_arith.v"
`include "./SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic.v"
`include "./SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff.v"
`include "./SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric.v"
`include "./SRC/lb/logical_tile_clb_mode_default__fle.v"
`include "./SRC/lb/logical_tile_clb_mode_clb_.v"
`include "./SRC/lb/logical_tile_mult_18_mode_default__mult_18_core_mode_mult_18x18__mult_18x18_slice_mode_default__mult_18x18.v"
`include "./SRC/lb/logical_tile_mult_18_mode_default__mult_18_core_mode_mult_18x18__mult_18x18_slice.v"
`include "./SRC/lb/logical_tile_mult_18_mode_default__mult_18_core.v"
`include "./SRC/lb/logical_tile_mult_18_mode_mult_18_.v"
// `include "./SRC/lb/grid_io_top_top.v"
// `include "./SRC/lb/grid_io_right_right.v"
// `include "./SRC/lb/grid_io_bottom_bottom.v"
// `include "./SRC/lb/grid_io_left_left.v"
`include "./SRC/lb/grid_clb.v"
`include "./SRC/lb/grid_mult_18.v"

// ------ Include routing module netlists -----
`include "./SRC/routing/sb_0__0_.v"
`include "./SRC/routing/sb_0__1_.v"
`include "./SRC/routing/sb_0__3_.v"
`include "./SRC/routing/sb_0__4_.v"
`include "./SRC/routing/sb_1__0_.v"
`include "./SRC/routing/sb_1__1_.v"
`include "./SRC/routing/sb_1__2_.v"
`include "./SRC/routing/sb_1__3_.v"
`include "./SRC/routing/sb_1__4_.v"
`include "./SRC/routing/sb_2__2_.v"
`include "./SRC/routing/sb_2__3_.v"
`include "./SRC/routing/sb_4__0_.v"
`include "./SRC/routing/sb_4__1_.v"
`include "./SRC/routing/sb_4__2_.v"
`include "./SRC/routing/sb_4__3_.v"
`include "./SRC/routing/sb_4__4_.v"
`include "./SRC/routing/cbx_1__0_.v"
`include "./SRC/routing/cbx_1__1_.v"
`include "./SRC/routing/cbx_1__4_.v"
`include "./SRC/routing/cbx_2__3_.v"
`include "./SRC/routing/cby_0__1_.v"
`include "./SRC/routing/cby_1__1_.v"
`include "./SRC/routing/cby_2__3_.v"
`include "./SRC/routing/cby_4__1_.v"
`include "./SRC/routing/cby_4__3_.v"

// ------ Include fabric top-level netlists -----
`include "./fpga_top_cocosim.v"

`include "./SRC/fpga_core.v"
//----- Include STD Cell netlists -----
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111o/sky130_fd_sc_hd__a2111o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2111oi/sky130_fd_sc_hd__a2111oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211o/sky130_fd_sc_hd__a211o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a211oi/sky130_fd_sc_hd__a211oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21bo/sky130_fd_sc_hd__a21bo_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21boi/sky130_fd_sc_hd__a21boi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21o/sky130_fd_sc_hd__a21o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a21oi/sky130_fd_sc_hd__a21oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221o/sky130_fd_sc_hd__a221o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a221oi/sky130_fd_sc_hd__a221oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a222oi/sky130_fd_sc_hd__a222oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a222oi/sky130_fd_sc_hd__a222oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a222oi/sky130_fd_sc_hd__a222oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a222oi/sky130_fd_sc_hd__a222oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22o/sky130_fd_sc_hd__a22o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a22oi/sky130_fd_sc_hd__a22oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2o/sky130_fd_sc_hd__a2bb2o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a2bb2oi/sky130_fd_sc_hd__a2bb2oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311o/sky130_fd_sc_hd__a311o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a311oi/sky130_fd_sc_hd__a311oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31o/sky130_fd_sc_hd__a31o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a31oi/sky130_fd_sc_hd__a31oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32o/sky130_fd_sc_hd__a32o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a32oi/sky130_fd_sc_hd__a32oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41o/sky130_fd_sc_hd__a41o_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/a41oi/sky130_fd_sc_hd__a41oi_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2/sky130_fd_sc_hd__and2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and2b/sky130_fd_sc_hd__and2b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3/sky130_fd_sc_hd__and3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and3b/sky130_fd_sc_hd__and3b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4/sky130_fd_sc_hd__and4_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4b/sky130_fd_sc_hd__and4b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/and4bb/sky130_fd_sc_hd__and4bb_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_12.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_6.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/buf/sky130_fd_sc_hd__buf_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufbuf/sky130_fd_sc_hd__bufbuf.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufbuf/sky130_fd_sc_hd__bufbuf.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufbuf/sky130_fd_sc_hd__bufbuf.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufbuf/sky130_fd_sc_hd__bufbuf_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufbuf/sky130_fd_sc_hd__bufbuf_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufinv/sky130_fd_sc_hd__bufinv.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufinv/sky130_fd_sc_hd__bufinv.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufinv/sky130_fd_sc_hd__bufinv.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufinv/sky130_fd_sc_hd__bufinv_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/bufinv/sky130_fd_sc_hd__bufinv_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkbuf/sky130_fd_sc_hd__clkbuf_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s15/sky130_fd_sc_hd__clkdlybuf4s15.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s15/sky130_fd_sc_hd__clkdlybuf4s15.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s15/sky130_fd_sc_hd__clkdlybuf4s15.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s15/sky130_fd_sc_hd__clkdlybuf4s15_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s15/sky130_fd_sc_hd__clkdlybuf4s15_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s18/sky130_fd_sc_hd__clkdlybuf4s18.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s18/sky130_fd_sc_hd__clkdlybuf4s18.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s18/sky130_fd_sc_hd__clkdlybuf4s18.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s18/sky130_fd_sc_hd__clkdlybuf4s18_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s18/sky130_fd_sc_hd__clkdlybuf4s18_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s25/sky130_fd_sc_hd__clkdlybuf4s25.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s25/sky130_fd_sc_hd__clkdlybuf4s25.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s25/sky130_fd_sc_hd__clkdlybuf4s25.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s25/sky130_fd_sc_hd__clkdlybuf4s25_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s25/sky130_fd_sc_hd__clkdlybuf4s25_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s50/sky130_fd_sc_hd__clkdlybuf4s50.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s50/sky130_fd_sc_hd__clkdlybuf4s50.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s50/sky130_fd_sc_hd__clkdlybuf4s50.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s50/sky130_fd_sc_hd__clkdlybuf4s50_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkdlybuf4s50/sky130_fd_sc_hd__clkdlybuf4s50_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinv/sky130_fd_sc_hd__clkinv_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinvlp/sky130_fd_sc_hd__clkinvlp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinvlp/sky130_fd_sc_hd__clkinvlp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinvlp/sky130_fd_sc_hd__clkinvlp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinvlp/sky130_fd_sc_hd__clkinvlp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/clkinvlp/sky130_fd_sc_hd__clkinvlp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/conb/sky130_fd_sc_hd__conb.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/conb/sky130_fd_sc_hd__conb.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/conb/sky130_fd_sc_hd__conb.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/conb/sky130_fd_sc_hd__conb_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap_12.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap_3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap_6.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/decap/sky130_fd_sc_hd__decap_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbn/sky130_fd_sc_hd__dfbbn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbn/sky130_fd_sc_hd__dfbbn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbn/sky130_fd_sc_hd__dfbbn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbn/sky130_fd_sc_hd__dfbbn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbn/sky130_fd_sc_hd__dfbbn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbp/sky130_fd_sc_hd__dfbbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbp/sky130_fd_sc_hd__dfbbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbp/sky130_fd_sc_hd__dfbbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfbbp/sky130_fd_sc_hd__dfbbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrbp/sky130_fd_sc_hd__dfrbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrbp/sky130_fd_sc_hd__dfrbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrbp/sky130_fd_sc_hd__dfrbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrbp/sky130_fd_sc_hd__dfrbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrbp/sky130_fd_sc_hd__dfrbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtn/sky130_fd_sc_hd__dfrtn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtn/sky130_fd_sc_hd__dfrtn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtn/sky130_fd_sc_hd__dfrtn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtn/sky130_fd_sc_hd__dfrtn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfrtp/sky130_fd_sc_hd__dfrtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfsbp/sky130_fd_sc_hd__dfsbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfsbp/sky130_fd_sc_hd__dfsbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfsbp/sky130_fd_sc_hd__dfsbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfsbp/sky130_fd_sc_hd__dfsbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfsbp/sky130_fd_sc_hd__dfsbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfstp/sky130_fd_sc_hd__dfstp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxbp/sky130_fd_sc_hd__dfxbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxbp/sky130_fd_sc_hd__dfxbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxbp/sky130_fd_sc_hd__dfxbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxbp/sky130_fd_sc_hd__dfxbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxbp/sky130_fd_sc_hd__dfxbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dfxtp/sky130_fd_sc_hd__dfxtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/diode/sky130_fd_sc_hd__diode.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/diode/sky130_fd_sc_hd__diode.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/diode/sky130_fd_sc_hd__diode.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/diode/sky130_fd_sc_hd__diode_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlclkp/sky130_fd_sc_hd__dlclkp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbn/sky130_fd_sc_hd__dlrbn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbn/sky130_fd_sc_hd__dlrbn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbn/sky130_fd_sc_hd__dlrbn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbn/sky130_fd_sc_hd__dlrbn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbn/sky130_fd_sc_hd__dlrbn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbp/sky130_fd_sc_hd__dlrbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbp/sky130_fd_sc_hd__dlrbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbp/sky130_fd_sc_hd__dlrbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbp/sky130_fd_sc_hd__dlrbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrbp/sky130_fd_sc_hd__dlrbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtn/sky130_fd_sc_hd__dlrtn_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlrtp/sky130_fd_sc_hd__dlrtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd1/sky130_fd_sc_hd__dlygate4sd1.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd1/sky130_fd_sc_hd__dlygate4sd1.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd1/sky130_fd_sc_hd__dlygate4sd1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd1/sky130_fd_sc_hd__dlygate4sd1_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd2/sky130_fd_sc_hd__dlygate4sd2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd2/sky130_fd_sc_hd__dlygate4sd2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd2/sky130_fd_sc_hd__dlygate4sd2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd2/sky130_fd_sc_hd__dlygate4sd2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd3/sky130_fd_sc_hd__dlygate4sd3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd3/sky130_fd_sc_hd__dlygate4sd3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd3/sky130_fd_sc_hd__dlygate4sd3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlygate4sd3/sky130_fd_sc_hd__dlygate4sd3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s2s/sky130_fd_sc_hd__dlymetal6s2s.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s2s/sky130_fd_sc_hd__dlymetal6s2s.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s2s/sky130_fd_sc_hd__dlymetal6s2s.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s2s/sky130_fd_sc_hd__dlymetal6s2s_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s4s/sky130_fd_sc_hd__dlymetal6s4s.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s4s/sky130_fd_sc_hd__dlymetal6s4s.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s4s/sky130_fd_sc_hd__dlymetal6s4s.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s4s/sky130_fd_sc_hd__dlymetal6s4s_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s6s/sky130_fd_sc_hd__dlymetal6s6s.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s6s/sky130_fd_sc_hd__dlymetal6s6s.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s6s/sky130_fd_sc_hd__dlymetal6s6s.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/dlymetal6s6s/sky130_fd_sc_hd__dlymetal6s6s_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ebufn/sky130_fd_sc_hd__ebufn_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxbp/sky130_fd_sc_hd__edfxbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxbp/sky130_fd_sc_hd__edfxbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxbp/sky130_fd_sc_hd__edfxbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxbp/sky130_fd_sc_hd__edfxbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxtp/sky130_fd_sc_hd__edfxtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxtp/sky130_fd_sc_hd__edfxtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxtp/sky130_fd_sc_hd__edfxtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/edfxtp/sky130_fd_sc_hd__edfxtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvn/sky130_fd_sc_hd__einvn_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/einvp/sky130_fd_sc_hd__einvp_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fa/sky130_fd_sc_hd__fa_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fah/sky130_fd_sc_hd__fah.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fah/sky130_fd_sc_hd__fah.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fah/sky130_fd_sc_hd__fah.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fah/sky130_fd_sc_hd__fah_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcin/sky130_fd_sc_hd__fahcin.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcin/sky130_fd_sc_hd__fahcin.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcin/sky130_fd_sc_hd__fahcin.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcin/sky130_fd_sc_hd__fahcin_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcon/sky130_fd_sc_hd__fahcon.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcon/sky130_fd_sc_hd__fahcon.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcon/sky130_fd_sc_hd__fahcon.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fahcon/sky130_fd_sc_hd__fahcon_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/fill/sky130_fd_sc_hd__fill_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/ha/sky130_fd_sc_hd__ha_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_12.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_6.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/inv/sky130_fd_sc_hd__inv_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_bleeder/sky130_fd_sc_hd__lpflow_bleeder.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_bleeder/sky130_fd_sc_hd__lpflow_bleeder.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_bleeder/sky130_fd_sc_hd__lpflow_bleeder.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_bleeder/sky130_fd_sc_hd__lpflow_bleeder_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkbufkapwr/sky130_fd_sc_hd__lpflow_clkbufkapwr_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_clkinvkapwr/sky130_fd_sc_hd__lpflow_clkinvkapwr_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr_12.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr_3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr_6.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_decapkapwr/sky130_fd_sc_hd__lpflow_decapkapwr_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0n/sky130_fd_sc_hd__lpflow_inputiso0n.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0n/sky130_fd_sc_hd__lpflow_inputiso0n.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0n/sky130_fd_sc_hd__lpflow_inputiso0n.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0n/sky130_fd_sc_hd__lpflow_inputiso0n_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0p/sky130_fd_sc_hd__lpflow_inputiso0p.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0p/sky130_fd_sc_hd__lpflow_inputiso0p.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0p/sky130_fd_sc_hd__lpflow_inputiso0p.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso0p/sky130_fd_sc_hd__lpflow_inputiso0p_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1n/sky130_fd_sc_hd__lpflow_inputiso1n.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1n/sky130_fd_sc_hd__lpflow_inputiso1n.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1n/sky130_fd_sc_hd__lpflow_inputiso1n.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1n/sky130_fd_sc_hd__lpflow_inputiso1n_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1p/sky130_fd_sc_hd__lpflow_inputiso1p.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1p/sky130_fd_sc_hd__lpflow_inputiso1p.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1p/sky130_fd_sc_hd__lpflow_inputiso1p.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputiso1p/sky130_fd_sc_hd__lpflow_inputiso1p_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputisolatch/sky130_fd_sc_hd__lpflow_inputisolatch.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputisolatch/sky130_fd_sc_hd__lpflow_inputisolatch.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputisolatch/sky130_fd_sc_hd__lpflow_inputisolatch.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_inputisolatch/sky130_fd_sc_hd__lpflow_inputisolatch_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrc/sky130_fd_sc_hd__lpflow_isobufsrc_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrckapwr/sky130_fd_sc_hd__lpflow_isobufsrckapwr.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrckapwr/sky130_fd_sc_hd__lpflow_isobufsrckapwr.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrckapwr/sky130_fd_sc_hd__lpflow_isobufsrckapwr.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/lpflow_isobufsrckapwr/sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/macro_sparecell/sky130_fd_sc_hd__macro_sparecell.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/macro_sparecell/sky130_fd_sc_hd__macro_sparecell.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/macro_sparecell/sky130_fd_sc_hd__macro_sparecell.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/maj3/sky130_fd_sc_hd__maj3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2/sky130_fd_sc_hd__mux2_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux2i/sky130_fd_sc_hd__mux2i_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/mux4/sky130_fd_sc_hd__mux4_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2/sky130_fd_sc_hd__nand2_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand2b/sky130_fd_sc_hd__nand2b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3/sky130_fd_sc_hd__nand3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand3b/sky130_fd_sc_hd__nand3b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4/sky130_fd_sc_hd__nand4_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4b/sky130_fd_sc_hd__nand4b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nand4bb/sky130_fd_sc_hd__nand4bb_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2/sky130_fd_sc_hd__nor2_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor2b/sky130_fd_sc_hd__nor2b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3/sky130_fd_sc_hd__nor3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor3b/sky130_fd_sc_hd__nor3b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4/sky130_fd_sc_hd__nor4_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4b/sky130_fd_sc_hd__nor4b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/nor4bb/sky130_fd_sc_hd__nor4bb_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111a/sky130_fd_sc_hd__o2111a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2111ai/sky130_fd_sc_hd__o2111ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211a/sky130_fd_sc_hd__o211a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o211ai/sky130_fd_sc_hd__o211ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21a/sky130_fd_sc_hd__o21a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ai/sky130_fd_sc_hd__o21ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21ba/sky130_fd_sc_hd__o21ba_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o21bai/sky130_fd_sc_hd__o21bai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221a/sky130_fd_sc_hd__o221a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o221ai/sky130_fd_sc_hd__o221ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22a/sky130_fd_sc_hd__o22a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o22ai/sky130_fd_sc_hd__o22ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2a/sky130_fd_sc_hd__o2bb2a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o2bb2ai/sky130_fd_sc_hd__o2bb2ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311a/sky130_fd_sc_hd__o311a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o311ai/sky130_fd_sc_hd__o311ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31a/sky130_fd_sc_hd__o31a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o31ai/sky130_fd_sc_hd__o31ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32a/sky130_fd_sc_hd__o32a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o32ai/sky130_fd_sc_hd__o32ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41a/sky130_fd_sc_hd__o41a_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/o41ai/sky130_fd_sc_hd__o41ai_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2_0.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2/sky130_fd_sc_hd__or2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or2b/sky130_fd_sc_hd__or2b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3/sky130_fd_sc_hd__or3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or3b/sky130_fd_sc_hd__or3b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4/sky130_fd_sc_hd__or4_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4b/sky130_fd_sc_hd__or4b_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/or4bb/sky130_fd_sc_hd__or4bb_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probec_p/sky130_fd_sc_hd__probec_p.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probec_p/sky130_fd_sc_hd__probec_p.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probec_p/sky130_fd_sc_hd__probec_p.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probec_p/sky130_fd_sc_hd__probec_p_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probe_p/sky130_fd_sc_hd__probe_p.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probe_p/sky130_fd_sc_hd__probe_p.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probe_p/sky130_fd_sc_hd__probe_p.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/probe_p/sky130_fd_sc_hd__probe_p_8.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbn/sky130_fd_sc_hd__sdfbbn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbn/sky130_fd_sc_hd__sdfbbn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbn/sky130_fd_sc_hd__sdfbbn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbn/sky130_fd_sc_hd__sdfbbn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbn/sky130_fd_sc_hd__sdfbbn_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbp/sky130_fd_sc_hd__sdfbbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbp/sky130_fd_sc_hd__sdfbbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbp/sky130_fd_sc_hd__sdfbbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfbbp/sky130_fd_sc_hd__sdfbbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrbp/sky130_fd_sc_hd__sdfrbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrbp/sky130_fd_sc_hd__sdfrbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrbp/sky130_fd_sc_hd__sdfrbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrbp/sky130_fd_sc_hd__sdfrbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrbp/sky130_fd_sc_hd__sdfrbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtn/sky130_fd_sc_hd__sdfrtn.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtn/sky130_fd_sc_hd__sdfrtn.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtn/sky130_fd_sc_hd__sdfrtn.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtn/sky130_fd_sc_hd__sdfrtn_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfrtp/sky130_fd_sc_hd__sdfrtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfsbp/sky130_fd_sc_hd__sdfsbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfsbp/sky130_fd_sc_hd__sdfsbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfsbp/sky130_fd_sc_hd__sdfsbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfsbp/sky130_fd_sc_hd__sdfsbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfsbp/sky130_fd_sc_hd__sdfsbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfstp/sky130_fd_sc_hd__sdfstp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxbp/sky130_fd_sc_hd__sdfxbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxbp/sky130_fd_sc_hd__sdfxbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxbp/sky130_fd_sc_hd__sdfxbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxbp/sky130_fd_sc_hd__sdfxbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxbp/sky130_fd_sc_hd__sdfxbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdfxtp/sky130_fd_sc_hd__sdfxtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sdlclkp/sky130_fd_sc_hd__sdlclkp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxbp/sky130_fd_sc_hd__sedfxbp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxbp/sky130_fd_sc_hd__sedfxbp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxbp/sky130_fd_sc_hd__sedfxbp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxbp/sky130_fd_sc_hd__sedfxbp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxbp/sky130_fd_sc_hd__sedfxbp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/sedfxtp/sky130_fd_sc_hd__sedfxtp_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor2/sky130_fd_sc_hd__xnor2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xnor3/sky130_fd_sc_hd__xnor3_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor2/sky130_fd_sc_hd__xor2_4.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3.behavioral.pp.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3.behavioral.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3_1.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3_2.v"
`include "/research/ece/lnis/CAD_TOOLS/DKITS/skywater/skywater-pdk/vendor/synopsys/PlaceRoute/sky130_fd_sc_hd/verilog/xor3/sky130_fd_sc_hd__xor3_4.v"
